    � B2SPICE zzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzz    ��  CPart          @           @                 74107D��  CIntPin    ��  CWire      �       �       �   �  p      �   �  p              74LS86N�    �    �   
   �         @           @                 74107D�    �    �      �         @           @                 74107D�    �    �       5  �        ��   TOutPort       _   @         _   @                 Output_Port ��  CExtPin    ��  CVertex3   �  `   ��  CSegment'    �-   �  `   �&   �   �  `                 �    �   �  `                                          �   port     �  �          Out1     ��   CPin                   ��                                                           @   port�� 
 TRectangle         �   `                   ����                                                 �   `   ��  TLine     @       @      ��       �                                                ��  TEllipse    8       H                  ����
[negative]               ���                       8       H      8       H   ��  
 TTextField (   ,   :   Q     ��                                                      (   ,   :   Q   (   ,   :   Q   [value]       �  $  0  �  (   ,   �   T   *�     $       <     ��                                                           $       <       $       <   [port.nbits]      <       ����            �      "Arial                    $       <   *�     ����j         ��                                                           ����j           ����j       	[refname]       �  �  �  (      �����       '   # ) + , - %      Output_Port     Miscellaneous      �?      ��   TOutPortModel       port ��  	 TModelPin ����port����        port����                                         0��    ��������             0��    ��������             0��    ��������             0��    ��������             0��    ��������             0��    �������� d   :�0�yE>10e-9��    �������� d   :�0�yE>10e-9��    ��������                             ����  ����:�0�yE>10e-9��d         ����  ����:�0�yE>10e-9��d   �      /   �����     ��   d   :�0�yE>10e-9��    �������� d   :�0�yE>10e-9��    ��������Output_PortOutput_Port   �            1 Digital<   Generic   Out1Out1           ����  ��    �������� ����  ��    �������� ����  ��    �������� ����  ��    �������� ����  ��    �������� ����  ��    �������� ����  ��    ��������  ��    ����       ����  Out ��   CPartPin    ����portport       A �      Digital Instruments Generic                                                                                                             5  1 0�    Q����   ����Q����                         �� �  :�0�ye>40ns��    ��������      x��    �������� �   I�����Z>25ns��    �������� �   I�����Z>25ns��    ��������      x��    �������� �   ��&�.Q>16ns��    �������� d   :�0�yE>10e-9��    �������� d   :�0�yE>10e-9��    ��������                            ����  ����:�0�yE>10e-9��d         ����  ����:�0�yE>10e-9��d   �      ��   TJKFF_general       JCkKRQQ' 0�     J����    ����J����                          ��      x��    ��������      x��    ��������      x��    ��������      x��    ��������      x��    ��������      x��    �������� d   :�0�yE>10e-9��    �������� d   :�0�yE>10e-9��    ��������                             ����  ����:�0�yE>10e-9��d         ����  ����:�0�yE>10e-9��d   �      6   �����     ��   d   :�0�yE>10e-9��    �������� d   :�0�yE>10e-9��    ��������0�    Ck����   ����Ck����                          ��      x��    ��������      x��    ��������      x��    ��������      x��    ��������      x��    ��������      x��    �������� d   :�0�yE>10e-9��    �������� d   :�0�yE>10e-9��    ��������                            ����  ����:�0�yE>10e-9��d         ����  ����:�0�yE>10e-9��d   �     �    �   9    11 �   9   �         @           @                 74107D�    
    < 13 ; �   �	    �   ?  	  14 >  0�    Q'����   ����Q'����                         �� �  :�0�ye>40ns��    ��������      x��    �������� �   I�����Z>25ns��    �������� �   I�����Z>25ns��    ��������      x��    �������� �   ��&�.Q>16ns��    �������� d   :�0�yE>10e-9��    �������� d   :�0�yE>10e-9��    ��������                           ����  ����:�0�yE>10e-9��d         ����  ����:�0�yE>10e-9��d   �     ? 5�       JCkKRQQ' 0�     J����    ����J����                          ��      x��    ��������      x��    ��������      x��    ��������      x��    ��������      x��    ��������      x��    �������� d   :�0�yE>10e-9��    �������� d   :�0�yE>10e-9��    ��������                             ����  ����:�0�yE>10e-9��d         ����  ����:�0�yE>10e-9��d   �      B   �����     ��   d   :�0�yE>10e-9��    �������� d   :�0�yE>10e-9��    ��������0�    Ck����   ����Ck����                          ��      x��    ��������      x��    ��������      x��    ��������      x��    ��������      x��    ��������      x��    �������� d   :�0�yE>10e-9��    �������� d   :�0�yE>10e-9��    ��������                            ����  ����:�0�yE>10e-9��d         ����  ����:�0�yE>10e-9��d   �     9 B   �����     ��   d   :�0�yE>10e-9��    �������� d   :�0�yE>10e-9��    ��������0�    K����   ����K����                          ��      x��    ��������      x��    ��������      x��    ��������      x��    ��������      x��    ��������      x��    �������� d   :�0�yE>10e-9��    �������� d   :�0�yE>10e-9��    ��������                             ����  ����:�0�yE>10e-9��d         ����  ����:�0�yE>10e-9��d   �     �    �   F    10 �   F    10  0�    Q'����   ����Q'����                         �� �  :�0�ye>40ns��    ��������      x��    �������� �   I�����Z>25ns��    �������� �   I�����Z>25ns��    ��������      x��    �������� �   ��&�.Q>16ns��    �������� d   :�0�yE>10e-9��    �������� d   :�0�yE>10e-9��    ��������                           ����  ����:�0�yE>10e-9��d         ����  ����:�0�yE>10e-9��d   �     F 5�       JCkKRQQ' 0�     J����    ����J����                          ��      x��    ��������      x��    ��������      x��    ��������      x��    ��������      x��    ��������      x��    �������� d   :�0�yE>10e-9��    �������� d   :�0�yE>10e-9��    ��������                             ����  ����:�0�yE>10e-9��d         ����  ����:�0�yE>10e-9��d   �      J   �����     ��   d   :�0�yE>10e-9��    �������� d   :�0�yE>10e-9��    ��������0�    Ck����   ����Ck����                          ��      x��    ��������      x��    ��������      x��    ��������      x��    ��������      x��    ��������      x��    �������� d   :�0�yE>10e-9��    �������� d   :�0�yE>10e-9��    ��������                            ����  ����:�0�yE>10e-9��d         ����  ����:�0�yE>10e-9��d   �     9 J   �����     ��   d   :�0�yE>10e-9��    �������� d   :�0�yE>10e-9��    ��������0�    K����   ����K����                          ��      x��    ��������      x��    ��������      x��    ��������      x��    ��������      x��    ��������      x��    �������� d   :�0�yE>10e-9��    �������� d   :�0�yE>10e-9��    ��������                             ����  ����:�0�yE>10e-9��d         ����  ����:�0�yE>10e-9��d   �     �    �   N    6 �   N    6  0�    Q'����   ����Q'����                         �� �  :�0�ye>40ns��    ��������      x��    �������� �   I�����Z>25ns��    �������� �   I�����Z>25ns��    ��������      x��    �������� �   ��&�.Q>16ns��    �������� d   :�0�yE>10e-9��    �������� d   :�0�yE>10e-9��    ��������                           ����  ����:�0�yE>10e-9��d         ����  ����:�0�yE>10e-9��d   �     N 6   �����        d   :�0�yE>10e-9��    �������� d   :�0�yE>10e-9��    ��������M  6J   �����     ��   d   :�0�yE>10e-9��    �������� d   :�0�yE>10e-9��    ��������0�    R����   ����R����                          ��      x��    ��������      x��    ��������      x��    ��������      x��    ��������      x��    ��������      x��    �������� d   :�0�yE>10e-9��    �������� d   :�0�yE>10e-9��    ��������                            ����  ����:�0�yE>10e-9��d         ����  ����:�0�yE>10e-9��d   �     �    �   S    12 �    S    ��   TInPort       _   @         _   @                 InputU �    �)   �   
   �    Y �6   �   
   �   �,   �  �   \         [     Z �   [ �    	   
   �   �+    	  �   `        _     ^ �   _ �	   `   
   �   �   `  �   d        c     �   c �   `   
   �   �*   `  �   h        g     f         b                                    @  �   A   �  `	          In1     "�                    ��                                                       �   @   A(� �   8   �   H                  ����
[negative]               ���                    �   8   �   H   �   8   �   H   $� t       �   @                   ����A                                      t       �   @   $� t   @   �   `                   ����A                                      t   @   �   `   &� �   @   �   @     ��                                                       $�         �   `                   ����                                                 �   `   &� t       t   `     
 ��                                                      ��  TPolygon                    ��                                                       ��  TPoint�   \    ��Ts��   P        s��   P       s��   D        s��   D        s��   P    ��Ks��   P    (�V    q�                    ��                                                       s��   $    hDWs��   0    �� s��   0    �  s��   <    �Qs��   <        s��   0    XKUs��   0    �OX    *� �       �   8    	 ��        	                                               �       �   8   �       �   8   	[A.nbits]      <       ����            �      "Arial                �       �   8   *�    (      M     ��        
                                                 (      M      (      M   [value]       �  �	  �  n
     (   l   P   *� ��������+   #     ��                                                       ��������+   #   ��������+   #   	[refname]       �  Q	  "  �	  ���������       j o   n   m {   � r � � l   k p ܕ    input_general     Miscellaneous      �?      ��   TInPortModel       A 0�     A����    ����A����                         ��             0��    ��������             0��    ��������             0��    ��������             0��    ��������             0��    ��������             0��    �������� d   :�0�yE>10e-9��    �������� d   :�0�yE>10e-9��    ��������                            ����  ����:�0�yE>10e-9��d         ����  ����:�0�yE>10e-9��d   �     S �   �����        d   :�0�yE>10e-9��    �������� d   :�0�yE>10e-9��    ��������1 Bit Inport1 Bit Inport   X            � Digital<   Generic   In1In1           ����  ��    �������� ����  ��    �������� ����  ��    �������� ����  ��    �������� ����  ��    �������� ����  ��    �������� ����  ��    ��������  X    ����            In 2�    ����AA      INAA�>  ����Digital Instruments Generic                         `   `              `   �  �              `   �             �  `   `          �      12 �   S    12 �   S    12 �   S   < 12  0�    R����   ����R����                          ��      x��    ��������      x��    ��������      x��    ��������      x��    ��������      x��    ��������      x��    �������� d   :�0�yE>10e-9��    �������� d   :�0�yE>10e-9��    ��������                            ����  ����:�0�yE>10e-9��d         ����  ����:�0�yE>10e-9��d   �     S 6   �����     ��   d   :�0�yE>10e-9��    �������� d   :�0�yE>10e-9��    ��������R 0�    R����   ����R����                          ��      x��    ��������      x��    ��������      x��    ��������      x��    ��������      x��    ��������      x��    �������� d   :�0�yE>10e-9��    �������� d   :�0�yE>10e-9��    ��������                            ����  ����:�0�yE>10e-9��d         ����  ����:�0�yE>10e-9��d   �     S B   �����     ��   d   :�0�yE>10e-9��    �������� d   :�0�yE>10e-9��    ��������0�    R����   ����R����                          ��      x��    ��������      x��    ��������      x��    ��������      x��    ��������      x��    ��������      x��    �������� d   :�0�yE>10e-9��    �������� d   :�0�yE>10e-9��    ��������                            ����  ����:�0�yE>10e-9��d         ����  ����:�0�yE>10e-9��d   �     S 5�       JCkKRQQ' 0�     J����    ����J����                          ��      x��    ��������      x��    ��������      x��    ��������      x��    ��������      x��    ��������      x��    �������� d   :�0�yE>10e-9��    �������� d   :�0�yE>10e-9��    ��������                             ����  ����:�0�yE>10e-9��d         ����  ����:�0�yE>10e-9��d   �     
 �   �����     ��   d   :�0�yE>10e-9��    �������� d   :�0�yE>10e-9��    ��������0�    Ck����   ����Ck����                          ��      x��    ��������      x��    ��������      x��    ��������      x��    ��������      x��    ��������      x��    �������� d   :�0�yE>10e-9��    �������� d   :�0�yE>10e-9��    ��������                            ����  ����:�0�yE>10e-9��d         ����  ����:�0�yE>10e-9��d   �     9 �   �����     ��   d   :�0�yE>10e-9��    �������� d   :�0�yE>10e-9��    ��������0�    K����   ����K����                          ��      x��    ��������      x��    ��������      x��    ��������      x��    ��������      x��    ��������      x��    �������� d   :�0�yE>10e-9��    �������� d   :�0�yE>10e-9��    ��������                             ����  ����:�0�yE>10e-9��d         ����  ����:�0�yE>10e-9��d   �     ? �   �����     ��   d   :�0�yE>10e-9��    �������� d   :�0�yE>10e-9��    ��������� 0�    Q����   ����Q����                         �� �  :�0�ye>40ns��    ��������      x��    �������� �   I�����Z>25ns��    �������� �   I�����Z>25ns��    ��������      x��    �������� �   ��&�.Q>16ns��    �������� d   :�0�yE>10e-9��    �������� d   :�0�yE>10e-9��    ��������                            ����  ����:�0�yE>10e-9��d         ����  ����:�0�yE>10e-9��d   �     �
    �   �  
 < 15 �    �   
 �       _   @         _   @                 Output_Port� �    �   @      �+   �0   @  �   �   �   �  `   �  
      �     �  
   �      
              �   port     @  @          Out4     "�                   ��                                                           @   port$�         �   `                   ����                                                 �   `   &�     @       @      ��                                                        (�    8       H                  ����
[negative]               ���                       8       H      8       H   *� (   ,   :   Q     ��                                                      (   ,   :   Q   (   ,   :   Q   [value]       �  �  �  Z  (   ,   �   T   *�     $       <     ��                                                           $       <       $       <   [port.nbits]      <       ����            �      "Arial                    $       <   *�     ����j         ��                                                           ����j           ����j       	[refname]       �  (  �  �      �����       �   � � � � � �      Output_Port     Miscellaneous      �?      .�       port 0� ����port����        port����                                         0��    ��������             0��    ��������             0��    ��������             0��    ��������             0��    ��������             0��    �������� d   :�0�yE>10e-9��    �������� d   :�0�yE>10e-9��    ��������                             ����  ����:�0�yE>10e-9��d         ����  ����:�0�yE>10e-9��d   �     � �   �����     ��   d   :�0�yE>10e-9��    �������� d   :�0�yE>10e-9��    ��������Output_PortOutput_Port   MJ            � Digital<   Generic   Out4Out4           ����  ��    �������� ����  ��    �������� ����  ��    �������� ����  ��    �������� ����  ��    �������� ����  ��    �������� ����  ��    ��������  10e-    ����       ����  Out 2�    ����portport       A �>      Digital Instruments Generic                                                                          -9��                                15  � � 
 15�   �����        d   :�0�yE>10e-9��    �������� d   :�0�yE>10e-9��    ��������0�    Q'����   ����Q'����                         �� �  :�0�ye>40ns��    ��������      x��    �������� �   I�����Z>25ns��    �������� �   I�����Z>25ns��    ��������      x��    �������� �   ��&�.Q>16ns��    �������� d   :�0�yE>10e-9��    �������� d   :�0�yE>10e-9��    ��������                           ����  ����:�0�yE>10e-9��d         ����  ����:�0�yE>10e-9��d   �     �    �   �   < 16 �   �    16  � 0� �  B����       B����                          ��      x��    ��������      x��    ��������      x��    ��������      x��    ��������      x��    ��������      x��    �������� d   :�0�yE>10e-9��    �������� d   :�0�yE>10e-9��    ��������                             ����  ����:�0�yE>10e-9��d         ����  ����:�0�yE>10e-9��d   �     � ��   TXOr       ABY 0� �  A����        A����                          ��      x��    ��������      x��    ��������      x��    ��������      x��    ��������      x��    ��������      x��    �������� d   :�0�yE>10e-9��    �������� d   :�0�yE>10e-9��    ��������                             ����  ����:�0�yE>10e-9��d         ����  ����:�0�yE>10e-9��d   �     
 �   �����     ��   d   :�0�yE>10e-9��    �������� d   :�0�yE>10e-9��    ��������� 0� �  Y����       Y����                         �� �   �U��T>19.5ns��    ��������      x��    �������� s   vԷ1�H>11.5ns��    �������� 	  gS��Ct\>26.5ns��    ��������      x��    �������� �   ��&�.Q>16ns��    �������� d   :�0�yE>10e-9��    �������� d   :�0�yE>10e-9��    ��������                            ����  ����:�0�yE>10e-9��d         ����  ����:�0�yE>10e-9��d   �      �   �����         d   :�0�yE>10e-9��    �������� d   :�0�yE>10e-9��    ��������86/4 LS 2-input XOr86/4 LS 2-input XOr   �            � � � Digital<   Generic   A6A6           ���� x��    �������� ���� x��    �������� � �h㈵�?40u��    �������� ��-C��6J�-.8m��    �������� ���,C��6:�-400u��    ��������  ������Mb�?8m��    �������� @ɢ�HP�x?6.1m��    ��������        ����LS      �����     ��   d   :�0�yE>10e-9��    �������� d   :�0�yE>10e-9��    �������� 16�   �����         d   :�0�yE>10e-9��    �������� d   :�0�yE>10e-9��    ��������107 JK FF w/clear107 JK FF w/clear                 � � � � � � Digital<   Generic   A4A4           ���� x��    �������� ���� x��    �������� �'	 hUMu?60u��    �������� ʑ�b2U0*�c�-2.4m��    �������� ���-C��6:�-.4m��    ��������  h�	����Mb�?16m��    ��������  ��{�G�z�?10m��    ��������  T��    ����Standard TTL                 0��    �������� ����    �sA20meg��    �������� 6  ��创�`>31n��    ��������             0��    ��������  �����     ��   d   :�0�yE>10e-9��    �������� d   :�0�yE>10e-9��    ���������  12J   �����     ��   d   :�0�yE>10e-9��    �������� d   :�0�yE>10e-9��    ��������0�    Q����   ����Q����                         �� �  :�0�ye>40ns��    ��������      x��    �������� �   I�����Z>25ns��    �������� �   I�����Z>25ns��    ��������      x��    �������� �   ��&�.Q>16ns��    �������� d   :�0�yE>10e-9��    �������� d   :�0�yE>10e-9��    ��������                            ����  ����:�0�yE>10e-9��d         ����  ����:�0�yE>10e-9��d   �      J   �����         d   :�0�yE>10e-9��    �������� d   :�0�yE>10e-9��    ��������I 107 JK FF w/clear107 JK FF w/clear                 K L M R � I Digital<   Generic   A2A2           ���� x��    �������� ���� x��    �������� �'	 hUMu?60u��    �������� ʑ�b2U0*�c�-2.4m��    �������� ���-C��6:�-.4m��    ��������  h�	����Mb�?16m��    ��������  ��{�G�z�?10m��    ��������  T��    ����Standard TTL                 0��    �������� ����    �sA20meg��    �������� 6  ��创�`>31n��    ��������             0��    ��������  �����        d   :�0�yE>10e-9��    �������� d   :�0�yE>10e-9��    ��������E  10B   �����     ��   d   :�0�yE>10e-9��    �������� d   :�0�yE>10e-9��    ��������� 0�    Q����   ����Q����                         �� �  :�0�ye>40ns��    ��������      x��    �������� �   I�����Z>25ns��    �������� �   I�����Z>25ns��    ��������      x��    �������� �   ��&�.Q>16ns��    �������� d   :�0�yE>10e-9��    �������� d   :�0�yE>10e-9��    ��������                            ����  ����:�0�yE>10e-9��d         ����  ����:�0�yE>10e-9��d   �     
 B   �����        d   :�0�yE>10e-9��    �������� d   :�0�yE>10e-9��    ��������A 107 JK FF w/clear107 JK FF w/clear                 C D E � � A Digital<   Generic   A3A3           ���� x��    �������� ���� x��    �������� �'	 hUMu?60u��    �������� ʑ�b2U0*�c�-2.4m��    �������� ���-C��6:�-.4m��    ��������  h�	����Mb�?16m��    ��������  ��{�G�z�?10m��    ��������  ��<     ����Standard TTL                 0��    �������� ����    �sA20meg��    �������� 6  ��创�`>31n��    ��������             0��    ��������  �����         d   :�0�yE>10e-9��    �������� d   :�0�yE>10e-9��    ��������� 	 14 	 < 14 � � � �    �   @  `   �"   �1   @      �    
     �     �   � �4   �  `   �   �   �  `   �        �     � �   � �9   �  �   �	   �   �  �   �     �     �                                    �  J�  �   �   @  �   �   �   �  �   �   �"   �  �   �     �     � �   � �    
  �   � �   � �&   @  �   �            �   � �   �  �   � �   � �'   �  �   �            �   � �      �   � �   �%   �  �   �         �     �   � �(   �  �   �                                         �                  �  Ck�  �   �   @      �#   �   �      �  	      �      	            @  K�  �   i         R�  �   �   @  �  Q�  �   �   �      �!   �          �     �     �   � �7   `      �(   �8   `      �*   �   �      �        �     �     �     �                  @  @  Q'�   @  �          A4     "�                    ��                                                           �   J"�                   ��                                                          �   Ck"�                   ��                                                          �   K"�                   ��                                                      `      R"�                   ��                                                      �   �   Q"�                   ��                                                      �   �   Q'$�     `   �   �                  ����                                             `   �   �   &�     �       �     ��       �                                                &�     �       �     ��                                                        &�     �       �    	 ��        	                                                &� `   �   `       
 ��       �
                                                &� �   �   �   �     ��                                                        &� �   �   �   �     ��                                                        &� �   x   �   �     ��                                                        &� �   x   �   x     ��                                                        (� X   �   h   �                  �                                           X   �   h   �   X   �   h   �   &� �   �   �   �     ��    ����                                                &� �   �   �   �     ��    ����                                                (� �   �   �   �                  �                                           �   �   �   �   �   �   �   �   *�     0   b   X     ��                                                           0   b   X       0   b   X   	[refname]       �  p  h        0   �   T   *� (   p   0   �     ��                                                      (   p   0   �   (   p   0   �   j       �  0  �  �  (   p   p   �   *� (   �   P   �     ��                                                      (   �   P   �   (   �   P   �   clk       �  �  0  &  (   �   p   �   *� (   �   8   �     ��                                                      (   �   8   �   (   �   8   �   k       �  �  �  �  (   �   p   �   *�        �   0     ��                                                              �   0          �   0   	[devname]        ����������������       �   0    � � � � � � � � � � � � � � � �       �   � � � � � �   �      74107 JK FF w/clear    74107 JK FF w/clear IEEEMiscellaneous      �?      �   A 2�    ����JJ      INAJ�C  ����2�   ����CkCk      INACk�C  ����2�   ����KK      INAK�C  ����2�   ����RR      INAR    ����2�   ����QQ      OUTAQT  ����2�   ����Q'Q'      OUTAQ'�>  ����2�    ����JJ      INBJ�>  ����2�   ����CkCk      INBCk�>  ����2�   ����KK      INBK�>  ����2�   ����RR      INBR�>  ����2�   ����QQ      OUTBQ�C  ����2�   ����Q'Q'      OUTBQ'�C  ����
Flip FlopsJK Flip-Flop w/clearGenericDO14             11 �   9    11 �   9    11 �    9    ��   TClock       �   �  �      �   �  �              Clock
�    �    �     A�      �          U2     "�                   ��                                                       �   `   A$�     @   �   �                  ����                                             @   �   �   &� �   `   �   `     ��                                                       &� `   @   `   �     ��    ����                                                &� p   h   x   h     ��                                                        &� x   T   x   h     ��       �                                                &� x   T   �   T     ��    ����                                                &� �   T   �   h     ��    ��T                                                &� �   h   �   h     ��    ��W                                                &� �   P   �   p      ��    ��W	                                                *�    P   Z   u    
 ��        
                                                  P   Z   u      P   Z   u   [period]       P  p  0  	     P   P   t   *� �   `   �   �    	 ��                                                      �   `   �   �   �   `   �   �   ns          �  p  6	  �   `   �   x   *�     �����        ��                                                           �����          �����      	[devname]        ����������������    �����      *�        *   @     ��                                                              *   @          *   @   	[refname]          �  �  h         �   <                             Clock     Miscellaneous      �?      ��   TClockModel     ��  CValue �  I�����z>100n      ��������� �  I�����j>50n     �������� A 0�     A����    ����A����                          ��      x��    ��������      x��    ��������      x��    ��������      x��    ��������      x��    ��������      x��    �������� d   :�0�yE>10e-9��    �������� d   :�0�yE>10e-9��    ��������                             ����  ����:�0�yE>10e-9��d         ����  ����:�0�yE>10e-9��d   �     9   �����         d   :�0�yE>10e-9��    �������� d   :�0�yE>10e-9��    ��������ClockClock   �          !Digital InstrumentsO   Generic   U2U2           ����  ��    �������� ����  ��    �������� ����  ��    �������� ����  ��    �������� ����  ��    �������� ����  ��    �������� ����  ��    ��������  `X    ����Generic             U 2�    ����AA      INAA    ����Digital InstrumentsDigital Clock inputGeneric                                                                                                                   11  8 L D � ! 116   �����     ��   d   :�0�yE>10e-9��    �������� d   :�0�yE>10e-9��    ��������0�    K����   ����K����                          ��      x��    ��������      x��    ��������      x��    ��������      x��    ��������      x��    ��������      x��    �������� d   :�0�yE>10e-9��    �������� d   :�0�yE>10e-9��    ��������                             ����  ����:�0�yE>10e-9��d         ����  ����:�0�yE>10e-9��d   �     �    �   $   3 �   $  �         �  �        �  �              7404D�         '1 &�    �   @      �   �!   �      +�
   �#   �  `   �   .�    �  `   /              �   �   �  �   �)   2�       �   3            1     .    -     ,         *                    �  in�  �   �$          �   6�   �      7                     �  �  out�   @  �          A5     "�                   ��                                                           �   in"�                   ��                                                      �   �   out(� l   t   �   �                   ���                                          l   t   �   �   l   t   �   �   &� �   �   �   �     ��                                                        &�     �   ,   �     ��    ����                                                q� ����    ����      ��                                                         s�,   \    XR�s�,   �       s�l   �    `  s�,   \     zW    *� ����   �   0     ��                                                       ����   �   0   ����   �   0   	[devname]        ��������������������   �   0   *� ����0   >   X     ��                                                       ����0   >   X   ����0   >   X   	[refname]       4  0  �  �  ����0   �   T   	 ;  9=:>CD<     Inverter    Inverter IEEEMiscellaneous      �?    =  ��   TAnd       InY 0�     In����    ����In����                          ��      x��    ��������      x��    ��������      x��    ��������      x��    ��������      x��    ��������      x��    �������� d   :�0�yE>10e-9��    �������� d   :�0�yE>10e-9��    ��������                             ����  ����:�0�yE>10e-9��d         ����  ����:�0�yE>10e-9��d   �      F  �����     ��   d   :�0�yE>10e-9��    �������� d   :�0�yE>10e-9��    ��������0�    Y����   ����Y����                         �� �   ,i�)+P>15ns��    ��������      x��    �������� d   :�0�yE>10ns��    �������� �   ,i�)+P>15ns��    ��������      x��    �������� Z   h�+e�SC>9ns��    �������� d   :�0�yE>10e-9��    �������� d   :�0�yE>10e-9��    ��������                           ����  ����:�0�yE>10e-9��d         ����  ����:�0�yE>10e-9��d   �     $F  �����        d   :�0�yE>10e-9��    �������� d   :�0�yE>10e-9��    ��������04/6 LS Inverter04/6 LS Inverter = �            GHDigital<   Generic   A5A5           ���� x��    �������� ���� x��    �������� @ �h㈵��>20u��    �������� ���-C��6:�-.4m��    �������� ���-C��6:�-.4m��    ��������  ������Mb�?8m��    ��������  6nb2U0*�c?2.4m��    ��������          ����LS      A 2�    ����inIn      PASA1A    ����2�   ����outY      PASA1Y   ����2�    ����inIn      PASB1A   ����2�   ����outY      PASB1Y   ����2�    ����inIn      PASC1A   ����2�   ����outY      PASC1Y   ����2�    ����inIn      PASD1A    ����2�   ����outY      PASD1Y   ����2�    ����inIn      PASE1A    ����2�   ����outY      PASE1Y0������2�    ����inIn      PASF1A  0����2�   ����outY      PASF1Y    ����Gatesdigital one-bit-wide inverterGenericDO14              3  #H 36   �����     ��   d   :�0�yE>10e-9��    �������� d   :�0�yE>10e-9��    ��������� 4 Q 107 JK FF w/clear107 JK FF w/clear                 7 8 #� 4 Q Digital<   Generic   A1A1           ���� x��    �������� ���� x��    �������� �'	 hUMu?60u��    �������� ʑ�b2U0*�c�-2.4m��    �������� ���-C��6:�-.4m��    ��������  h�	����Mb�?16m��    ��������  ��{�G�z�?10m��    ��������  ��t    ����Standard TTL                 0��    �������� ����    �sA20meg��    �������� 6  ��创�`>31n��    ��������             0��    ��������  �����         d   :�0�yE>10e-9��    �������� d   :�0�yE>10e-9��    ��������K  5    5 	P �  G �            �  J�  �   �       �  Ck�  �   �   �      �   �   �      Y        X                 @  K�  �   a         R�  �   �    
  `   �   ]�.   �
  `   �$   �   @  `   `        _    ^�%   �2   �
  `   b   	     _                     @  �  Q�  �   �
    
      �   e�   @      f                    @  @  Q'�   �  �          A2     "�                    ��                                                           �   J"�                   ��                                                          �   Ck"�                   ��                                                          �   K"�                   ��                                                      `      R"�                   ��                                                      �   �   Q"�                   ��                                                      �   �   Q'$�     `   �   �                  ����                                             `   �   �   &�     �       �     ��                                                        &�     �       �     ��                                                        &�     �       �    	 ��        	                                                &� `   �   `       
 ��        
                                                &� �   �   �   �     ��                                                        &� �   �   �   �     ��                                                        &� �   x   �   �     ��                                                        &� �   x   �   x     ��                                                        (� X   �   h   �                  �                                           X   �   h   �   X   �   h   �   &� �   �   �   �     ��                                                        &� �   �   �   �     ��                                                        (� �   �   �   �                  �                                           �   �   �   �   �   �   �   �   *�     0   b   X     ��                                                           0   b   X       0   b   X   	[refname]       @  p  	        0   �   T   *� (   p   0   �     ��                                                      (   p   0   �   (   p   0   �   j       X  0  p  �  (   p   p   �   *� (   �   P   �     ��                                                      (   �   P   �   (   �   P   �   clk       X  �  �  &  (   �   p   �   *� (   �   8   �     ��                                                      (   �   8   �   (   �   8   �   k       X  �  �  �  (   �   p   �   *�        �   0     ��                                                              �   0          �   0   	[devname]        ����������������       �   0    hijklmnopqrst|}~      v  xyuz{  w     74107 JK FF w/clear    74107 JK FF w/clear IEEEMiscellaneous      �?      J   A 2�    ����JJ      INAJ�C  ����2�   ����CkCk      INACk��������2�   ����KK      INAK�C  ����2�   ����RR      INAR��������2�   ����QQ      OUTAQ   ����2�   ����Q'Q'      OUTAQ'   ����2�    ����JJ      INBJ�� �����2�   ����CkCk      INBCk��������2�   ����KK      INBKrier����2�   ����RR      INBRrial����2�   ����QQ      OUTBQ  � ����2�   ����Q'Q'      OUTBQ'   ����
Flip FlopsJK Flip-Flop w/clearGenericDO14             9  �        �	       _   @         _   @                 Output_Port��    c       �   port     �
  �          Out2     "�                   ��                                                           @   port$�         �   `                   ����                                                 �   `   &�     @       @      ��    `                                                   (�    8       H                  ����
[negative]               ���                       8       H      8       H   *� (   ,   :   Q     ��                                                      (   ,   :   Q   (   ,   :   Q   [value]       �
  $  0  �  (   ,   �   T   *�     $       <     ��                                                           $       <       $       <   [port.nbits]      <       ����            �      "Arial                    $       <   *�     ����j         ��                                                           ����j           ����j       	[refname]       �
  �  �  (      �����       �  ������     Output_Port     Miscellaneous      �?      .�       port 0� ����port����        port����                                         0��    ��������             0��    ��������             0��    ��������             0��    ��������             0��    ��������             0��    �������� d   :�0�yE>10e-9��    �������� d   :�0�yE>10e-9��    ��������                             ����  ����:�0�yE>10e-9��d         ����  ����:�0�yE>10e-9��d   �      �  �����     ��   d   :�0�yE>10e-9��    �������� d   :�0�yE>10e-9��    ��������Output_PortOutput_Port   MJ            �Digital<   Generic   Out2Out2           ����  ��    �������� ����  ��    �������� ����  ��    �������� ����  ��    �������� ����  ��    �������� ����  ��    �������� ����  ��    ��������          ����       ����  Out 2�    ����portport       A V      Digital Instruments Generic                                                                                                             9  �� C  9    9 H �  @ �    a       �  J�  �   �       �  Ck�  �   g      @  K�  �   e         R�  �   �   @  �  Q�  �   �   @  @  Q'�   @  �          A3     "�                    ��                                                           �   J"�                   ��                                                          �   Ck"�                   ��                                                          �   K"�                   ��                                                      `      R"�                   ��                                                      �   �   Q"�                   ��                                                      �   �   Q'$�     `   �   �                  ����                                             `   �   �   &�     �       �     ��                                                        &�     �       �     ��    �U                                                &�     �       �    	 ��    ���	                                                &� `   �   `       
 ��    �/ �
                                                &� �   �   �   �     ��                                                        &� �   �   �   �     ��                                                        &� �   x   �   �     ��     
 C                                                &� �   x   �   x     ��    P �                                                (� X   �   h   �                  �                                           X   �   h   �   X   �   h   �   &� �   �   �   �     ��     ���                                                &� �   �   �   �     ��    ���]                                                (� �   �   �   �                  �                                           �   �   �   �   �   �   �   �   *�     0   b   X     ��                                                           0   b   X       0   b   X   	[refname]       �  p  h        0   �   T   *� (   p   0   �     ��                                                      (   p   0   �   (   p   0   �   j       �  0  �  �  (   p   p   �   *� (   �   P   �     ��                                                      (   �   P   �   (   �   P   �   clk       �  �  0  &  (   �   p   �   *� (   �   8   �     ��                                                      (   �   8   �   (   �   8   �   k       �  �  �  �  (   �   p   �   *�        �   0     ��                                                              �   0          �   0   	[devname]        ����������������       �   0    ����������������      �  ������  �     74107 JK FF w/clear    74107 JK FF w/clear IEEEMiscellaneous      �?      B   A 2�    ����JJ      INAJ@  ����2�   ����CkCk      INACk    ����2�   ����KK      INAKAri����2�   ����RR      INAR    ����2�   ����QQ      OUTAQ�C  ����2�   ����Q'Q'      OUTAQ'�C  ����2�    ����JJ      INBJ�C  ����2�   ����CkCk      INBCk�C  ����2�   ����KK      INBK�C  ����2�   ����RR      INBR    ����2�   ����QQ      OUTBQ    ����2�   ����Q'Q'      OUTBQ'    ����
Flip FlopsJK Flip-Flop w/clearGenericDO14              13 = 	 �    
    �
       _   @         _   @                 Output_Port��    �        �   port     @  @          Out3     "�                   ��                                                           @   port$�         �   `                   ����                                                 �   `   &�     @       @      ��                                                       (�    8       H                  ����
[negative]               ���                       8       H      8       H   *� (   ,   :   Q     ��                                                      (   ,   :   Q   (   ,   :   Q   [value]       �  �  �  Z  (   ,   �   T   *�     $       <     ��                                                           $       <       $       <   [port.nbits]      <       ����            �      "Arial                    $       <   *�     ����j         ��                                                           ����j           ����j       	[refname]       �  (  �  �      �����       �  ������     Output_Port     Miscellaneous      �?      .�       port 0� ����port����        port����                                         0��    ��������             0��    ��������             0��    ��������             0��    ��������             0��    ��������             0��    �������� d   :�0�yE>10e-9��    �������� d   :�0�yE>10e-9��    ��������                             ����  ����:�0�yE>10e-9��d         ����  ����:�0�yE>10e-9��d   �     
 �  �����     ��   d   :�0�yE>10e-9��    �������� d   :�0�yE>10e-9��    ��������Output_PortOutput_Port   MJ            �Digital<   Generic   Out3Out3           ����  ��    �������� ����  ��    �������� ����  ��    �������� ����  ��    �������� ����  ��    �������� ����  ��    �������� ����  ��    ��������          ����       ����  Out 2�    ����portport       A V      Digital Instruments Generic                                                                                                             13  �� � �  13    13 �  �    �    �  �  a    �   �   �     b   �   4      �  y                 A6     "�                   ��                                                       �   �   a"�                   ��                                                      �   `   b"�                    ��                                                          �   y��   TArc ����p   d   �    	                                                              P   �   �      P   �   �   \   P      �           &� �   �   \   �     ��                                                        ց �����   d                                                                    0   �   �      0   �   �      �   \   �           &� �   P   \   P     ��                                                        &�     �       �     ��                                                        &� �   �   t   �     ��    e va                                                &� �   `   t   `     ��        	                                                ց �����      �    
           
                                                p   P   �   �   p   P   �   �   |   P   |   �           ց �����      �                                                               |   P   �   �   |   P   �   �   �   P   �   �           *�         �   (     ��                                                               �   (           �   (   	[devname]        ����������������        �   (   *�     $   B   L     ��                                                           $   B   L       $   B   L   	[refname]          l  �        $   �   H    �  ����  �  �����  �  �  �   XOR 2    
XOR 2 IEEEMiscellaneous      �?      �   A 2�    ����aA      INA1AT      2�   ����bB      INA1BU     2�   ����yY      OUTA1Y       2�    ����aA      INB1A        2�   ����bB      INB1B       2�   ����yY      OUTB1Y       2�    ����aA      INC1A        2�   ����bB      INC1BU     2�   ����yY      OUTC1YT     2�    ����aA      IND1AV      2�   ����bB      IND1B       2�   ����yY      OUTD1Y   �   Gatesquad 2-input xor gatesGenericDIP-14              1 ( 7 G�   1  �� 1 : %T  O �    0       �  J�  �   �       �  Ck�  �   8      @  K�  �   ]         R�  �   !   @  �  Q�  �   Z  @  @  Q'�   �  �          A1     "�                    ��                                                           �   J"�                   ��                                                          �   Ck"�                   ��                                                          �   K"�                   ��                                                      `      R"�                   ��                                                      �   �   Q"�                   ��                                                      �   �   Q'$�     `   �   �                  ����                                             `   �   �   &�     �       �     ��    �0S                                                &�     �       �     ��    @��                                                &�     �       �    	 ��    �7S	                                                &� `   �   `       
 ��    ��
                                                &� �   �   �   �     ��    P                                                  &� �   �   �   �     ��    �                                                &� �   x   �   �     ��    d                                                  &� �   x   �   x     ��    �a �                                                (� X   �   h   �                  �                                           X   �   h   �   X   �   h   �   &� �   �   �   �     ��    x                                                  &� �   �   �   �     ��    �1S                                                (� �   �   �   �                  �                                           �   �   �   �   �   �   �   �   *�     0   b   X     ��                                                           0   b   X       0   b   X   	[refname]       �  p  �        0   �   T   *� (   p   0   �     ��                                                      (   p   0   �   (   p   0   �   j       �  0    �  (   p   p   �   *� (   �   P   �     ��                                                      (   �   P   �   (   �   P   �   clk       �  �  p  &  (   �   p   �   *� (   �   8   �     ��                                                      (   �   8   �   (   �   8   �   k       �  �  (  �  (   �   p   �   *�        �   0     ��                                                              �   0          �   0   	[devname]        ����������������       �   0    ������������ 	
          0     74107 JK FF w/clear    74107 JK FF w/clear IEEEMiscellaneous      �?      6   A 2�    ����JJ      INAJU  ����2�   ����CkCk      INACk�  ����2�   ����KK      INAK0������2�   ����RR      INARB�r����2�   ����QQ      OUTAQ    ����2�   ����Q'Q'      OUTAQ'U  ����2�    ����JJ      INBJT  ����2�   ����CkCk      INBCk    ����2�   ����KK      INBK    ����2�   ����RR      INBR    ����2�   ����QQ      OUTBQX��K����2�   ����Q'Q'      OUTBQ'� �r����
Flip FlopsJK Flip-Flop w/clearGenericDO14                <   W ' ���      9 $S  N  F 
 ? � � , + ,   Y^f  � � � � � -1+� /7� � � � � � � � � \ h b ` f d ^ Z � � � `b  � 3� � : 7 : 0� 8� Z] � Xc eg a� g_ � � � � � e �   2� � ! � � *� 4,� .6� � � � Y i a ]  _  � � c �   [ � � �              
 �@ ����        ���������             0     ��������� ����      @5     ���������  ʚ;�������?.1     ���������@ ����       ��������� ����       ��������� ����       ��������� ����       ��������� ���� true
     ��������� ����  false     ��������               
                  � ����        ��������� ����       ���������  ����       ���������@ ����       ���������@ ����       ��������               
                  � ����        ��������� ����       ���������@ ����       ���������  ����       ��������� ����       ��������� ����       ��������� ����       ��������� ����       ��������� ����       ��������� ����       ��������� ����       ��������               
                 � ����dec     ��������� ����     @�@1k     ��������� ����    ��.A1meg     ��������� ����       20     ��������� ���� true     ��������� ���� true     ��������� ���� true	     ��������� ����  false
     ��������               
                 �  ����        ���������  ����       ���������  ����       ��������� ����dec     ��������� ����       ��������� ����       ��������� ����  	     ��������� ����  
     ��������               
                  	 � ����        ��������� ����       ��������� ����       ��������� ����       ��������� ����       ��������� ����       ��������� ����       ��������� ����       ��������� ����       ��������               
                 � ����        ��������� ����       ��������� ����       ��������� ����dec     ��������� ����       ��������               
                    �             0      ��������� ��� ����MbP?1m     ��������� �� �h㈵��>10u     ��������� '  ���ư>1u     ��������� ���� true     ��������� ����  false     ��������� ���� true     ��������� ����  false     ��������               
                 � ����     @�@1K      ���������  ����       ���������  ����       ���������  ����       ��������               
         ��              �  ����        ��������              
                  �  ����        ��������              
                                  
                 �@ ����        ���������@ ����       ��������� ����       ��������� ����       ��������� ����       ��������� ����       ��������� ����       ��������� ����       ��������� ����       ��������� ���� true	     ��������� ����  false
     ��������� ���� true     ��������� ����  false     ��������               
                 � ����       5      ��������� ����       5     ��������� ����       5     ��������� ����       5     ��������� ����       ��������� ����  	     ��������� ����  
     ��������� ����       ��������� ����       ��������� ����       ��������� ���� true     ���������@ ����       ���������@ ����       ��������� ����       ��������� ����       ��������� ����       ��������� ����dec     ��������� ����       ��������� ����       ��������� ����       ��������� ���� true     ��������� ���� true     ��������� ���� true     ��������� ����  false     ��������� ���� true     ��������� ����  false      ��������� ���� true!     ��������� ����  false"     ��������               
                        � ����       5      ��������� ����       5     ��������� ����       5     ��������� ����       5     ��������� ����       ��������� ����  	     ��������� ����  
     ��������� ����       ��������� ����       ��������� ����       ��������� ���� true     ���������@ ����       ���������@ ����       ��������� ����       ��������� ����       ��������� ����       ��������� ����dec     ��������� ����       ��������� ����       ��������� ����       ��������� ���� true     ��������� ���� true     ��������� ���� true     ��������� ����  false     ��������� ���� true     ��������� ����  false      ��������� ���� true!     ��������� ����  false"     ��������               
                 � ����       5      ��������� ����       5     ��������� ����       5     ��������� ����       5     ��������� ����       ��������� ����  	     ��������� ����  
     ��������� ����       ��������� ����       ��������� ����       ��������� ���� true     ���������@ ����       ���������@ ����       ��������� ����       ��������� ����       ��������� ����       ��������� ����dec     ��������� ����       ��������� ����       ��������� ����       ��������� ���� true     ��������� ���� true     ��������� ���� true     ��������� ����  false     ��������� ���� true     ��������� ����  false      ��������� ���� true!     ��������� ����  false"     ��������               
                 � ����       5      ��������� ����       5     ��������� ����       5     ��������� ����       5     ��������� ����       ��������� ����  	     ��������� ����  
     ��������� ����       ��������� ����       ��������� ����       ��������� ���� true     ���������@ ����       ���������@ ����       ��������� ����       ��������� ����       ��������� ����       ��������� ����dec     ��������� ����       ��������� ����       ��������� ����       ��������� ���� true     ��������� ���� true     ��������� ���� true     ��������� ����  false     ��������� ���� true     ��������� ����  false      ��������� ���� true!     ��������� ����  false"     ��������               
                 �@ ����        ���������@ ����       ��������� ����       ��������� ����       ��������� ����       ��������� ����       ��������� ����       ��������� ����       ��������� ����decade     ��������� ���� true     ��������� ���� true     ��������� ���� true     ��������� ����  false     ��������               
                 � ����        ��������� ����       ���������@ ����       ���������  ����       ��������� ����       ��������� ����       ��������� ����       ��������� ����       ��������� ����       ��������� ����       ��������� ����       ��������               
                        � ����dec     ��������� ����     @�@1k     ��������� ����    ��.A1meg     ��������� ����       20     ��������� ����        0     ��������� ����        0     ��������� ���� true	     ��������� ���� true
     ��������� ����      I@50     ��������� ���� true     ��������� ����  false     ��������               
                          / � ���� x'     ���������     �-���q=1E-12     ��������� @B -C��6?1E-4     ��������� ���� x     ��������� ���� x     ��������� ���� x     ��������� ���� x     ��������� ���� x     ��������� ���� x     ��������� ���� x	     ��������� ���� x!     ��������� ����    �  500
     ��������� ���� x     ��������� ����    �  500     ��������� ���� x$     ��������� ���� x$     ��������� ���� x%     ��������� ���� x"     ���������  ���� x*     ��������� ���� x     ��������� ���� x     ��������� ���� x     ��������� ���� x&     ��������� ���� x     ��������� ���� x     ��������� ���� x     ��������� ���� x+     ��������� ���� x,     ��������� ���� x-     ��������� ���� xg     ��������� ���� xf     ��������� ���� xd     ��������� ���� xe     ��������� ���� xh     ��������� ���� xj     ��������� ���� xi     ��������� ���� xk     ��������� ����    e��A1Gl     ���������             0�     ��������� ����      @5�     ��������� ����      @2.5�     ��������� ����      �?.5�     ��������� ����      @4.5�     ��������� 
   ��&�.>1n�     ��������� 
   ��&�.>1n�     ��������� 
   ��&�.>1n�     ��������� 
   ��&�.>1n�     ��������                                  Ariald        �ڬt�3Zx�  ۬t,� ���t    �ڬt�3Zx�  ۬t,� ���t ��  COpAnal                         
                        ����                                   �ڬt�3Zx�  ۬t,� ���t    �ڬt�3Zx�  ۬t,� ���t ��  CDCsweep       
  !               
                      ����                                   �ڬt�3Zx�  ۬t,� ���t    �ڬt�3Zx�  ۬t,� ���t ��  CACsweep        23456789               
                      ����                                  �ڬt�3Zx�  ۬t,� ���t    �ڬt�3Zx�  ۬t,� ���t �� 
 CTranSweep        PQRSTUVW               
                      ����                                   �ڬt�3Zx�  ۬t,� ���t    �ڬt�3Zx�  ۬t,� ���t ��  CACdisto        KLMNO               
                         ����                                  �ڬt�3Zx�  ۬t,� ���t    �ڬt�3Zx�  ۬t,� ���t 5�        � ����        ��������� ����       ��������� ����       ��������� ����dec     ��������� ����       ��������               
                          ����                                  �ڬt�3Zx�  ۬t,� ���t    �ڬt�3Zx�  ۬t,� ���t 5�        � ����        ��������� ����       ��������� ����       ��������� ����dec     ��������� ����       ��������               
                          ����                                  �ڬt�3Zx�  ۬t,� ���t    �ڬt�3Zx�  ۬t,� ���t 5�        � ����        ��������� ����       ��������� ����       ��������� ����dec     ��������� ����       ��������               
                          ����                                  �ڬt�3Zx�  ۬t,� ���t    �ڬt�3Zx�  ۬t,� ���t 5�        � ����        ��������� ����       ��������� ����       ��������� ����dec     ��������� ����       ��������               
                          ����                                  �ڬt�3Zx�  ۬t,� ���t    �ڬt�3Zx�  ۬t,� ���t 5�        � ����        ��������� ����       ��������� ����       ��������� ����dec     ��������� ����       ��������               
         �            	    ����                                  �ڬt�3Zx�  ۬t,� ���t    �ڬt�3Zx�  ۬t,� ���t ��  CACnoise        :;<=>?@A               
                   
    ����                                  �ڬt�3Zx�  ۬t,� ���t    �ڬt�3Zx�  ۬t,� ���t U�         �  ����        ���������  ����       ���������  ����       ��������� ����dec     ��������� ����       ��������� ����       ��������� ����  	     ��������� ����  
     ��������              
                        ����                                  �ڬt�3Zx�  ۬t,� ���t    �ڬt�3Zx�  ۬t,� ���t ��  CFourier        XYZ[               
         ��                  ����                                  �ڬt�3Zx�  ۬t,� ���t    �ڬt�3Zx�  ۬t,� ���t ��  CACpz        	 BCDEFGHIJ               
                       ����                                   �ڬt�3Zx�  ۬t,� ���t    �ڬt�3Zx�  ۬t,� ���t ��  CDCtf         "#$%&               
                       ����                                   �ڬt�3Zx�  ۬t,� ���t    �ڬt�3Zx�  ۬t,� ���t ��  CDCsens         '()*+,-./01               
                       ����                                   �ڬt�3Zx�  ۬t,� ���t    �ڬt�3Zx�  ۬t,� ���t                 ����                                  �ڬt�3Zx�  ۬t,� ���t    �ڬt�3Zx�  ۬t,� ���t ��  CShow         \              
                       ����                                   �ڬt�3Zx�  ۬t,� ���t    �ڬt�3Zx�  ۬t,� ���t ��  CShowmod         ]              
                       ����              0                   �ڬt�3Zx�  ۬t,� ���t    �ڬt�3Zx�  ۬t,� ���t �� 
 CLinearize        �  ����        ��������               
                      ����            �t�                   �ڬt�3Zx�  ۬t,� ���t    �ڬt�3Zx�  ۬t,� ���t ��  CParamTranSweep        ^_`abcdefghij               
                      ����             0�                   �ڬt�3Zx�  ۬t,� ���t    �ڬt�3Zx�  ۬t,� ���t 0             ����             2                     �ڬt�3Zx�  ۬t,� ���t    �ڬt�3Zx�  ۬t,� ���t ��  CParamACSweep        �������������               
                      ����                                  �ڬt�3Zx�  ۬t,� ���t    �ڬt�3Zx�  ۬t,� ���t ��  CMonteCarlo_op        klmnopqrstuvwxyz{|}~�������               
                             ����                                  �ڬt�3Zx�  ۬t,� ���t    �ڬt�3Zx�  ۬t,� ���t ��  CMonteCarlo_dc        ����������������������������               
                      ����                                   �ڬt�3Zx�  ۬t,� ���t    �ڬt�3Zx�  ۬t,� ���t ��  CMonteCarlo_ac        ����������������������������               
                      ����                                  �ڬt�3Zx�  ۬t,� ���t    �ڬt�3Zx�  ۬t,� ���t ��  CMonteCarlo_tran        ����������������������������               
                      ����                                   �ڬt�3Zx�  ۬t,� ���t    �ڬt�3Zx�  ۬t,� ���t ��  CACsens        �����������               
                             ����                                  �ڬt�3Zx�  ۬t,� ���t    �ڬt�3Zx�  ۬t,� ���t ��  CNetworkAnalysis        �����������               
                      ����                                  �ڬt�3Zx�  ۬t,� ���t    �ڬt�3Zx�  ۬t,� ���t                 ����                                >           ��   CDigSimResTemplate                 ��   TDigitalSignal            In1    ���� ����                        ��            U2    ���� ����                        ��            Out1    ���� ����                        ��            Out2    ���� ����                        ��            Out3    ���� ����                        ��            Out4    ���� ����                                 ���       ����  ����:�0�yU>+20.00n���   ����                       Arial����                       Arial����                       Arial                                           ����  ���� ������       ����  ���� ������                 �               ����  �����       200������          0.000000e+000��    ��������      0.000000e+000��    ��������      0.000000e+000��    ��������   ����                       Arial����                       Arial����                       Arial����                       Arial                        �     �   �  �                     ����  ��    ��������   @  DO14�14 pin small outline package                                                                                                                                                                                                                              ����   ��   CPackageAliasSuperPCBStandardSO14      ��EagleBURR.LBRSO14      ��Orcad SOG.050/14/WG.244/L.350      ��Pads SO14NB      ��	UltiboardL7IC.l55$SO14      ��Eagleburr-brown.lbrSO14             A              @  DO14�14 pin small outline package                                                                                                                                                                                                                              ����   ������        B              @  DO14�14 pin small outline package                                                                                                                                                                                                                              ����   ��SuperPCBStandardSO14      ��EagleBURR.LBRSO14      ��Orcad SOG.050/14/WG.244/L.350      ��Pads SO14NB      ��	UltiboardL7IC.l55$SO14      ��Eagleburr-brown.lbrSO14             A              @  DO14�14 pin small outline package                                                                                                                                                                                                                              ����   ������        B                                      @  DO14�14 pin small outline package                                                                                                                                                                                                                              ����   ��SuperPCBStandardSO14      ��EagleBURR.LBRSO14      ��Orcad SOG.050/14/WG.244/L.350      ��Pads SO14NB      ��	UltiboardL7IC.l55$SO14      ��Eagleburr-brown.lbrSO14             A                                                      �   DIP-14�14 pin dual in line package                                                                                                                                                                                                                               �     ��SuperPCBStandardDIP14      ��EagleBURR.LBRDIP-14      ��Orcad DIP.100/14/W.300/L.700      ��Pads DIP14      ��	UltiboardUltilib.l55DIP14      ��Eagleburr-brown.lbrDIL14      ��Eagledil.lbrDIL14     ��Eagleanalog-devicesDIL14      ��Eagle74xx-usDIL14      ��Eagle	74ttl-dinDIL14      ��EaglemaximDIL14      ��EagleexarDIL14      ��Eagle
ic-packageDIL14      ��Eagleresistor-dilDIL14      ��EagletexasDIL14      ��Eagle
74ac-logicDIL14              A      �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                   �#     ����t� xa	    <�     J   J   ��     xa	J                  2         �                 � � �           u m     ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                   �#     ����t� xa	    <�     J   J   ��     xa	J                  2         �                 � � �           u m     ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                   �#     ����t� xa	    <�     J   J   ��     xa	J                  2         �                 � � �           u m     ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                   �#     ����t� xa	    <�     J   J   ��     xa	J                  2         �                 � � �           u m     ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                   �#     ����t� xa	    <�     J   J   ��     xa	J                  2         �                 � � �           u m     ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                   �#     ����t� xa	    <�     J   J   ��     xa	J                  2         �                 � � �           u m     ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                   �#     ����t� xa	    <�     J   J   ��     xa	J                  2         �                 � � �           u m     ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                   �#     ����t� xa	    <�     J   J   ��     xa	J                  2         �                 � � �           u m     ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                   �#     ����t� xa	    <�     J   J   ��     xa	J                  2         �                 � � �           u m     ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                   �#     ����t� xa	    <�     J   J   ��     xa	J                  2         �                 � � �           u m     ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                   �#     ����t� xa	    <�     J   J   ��     xa	J                  2         �                 � � �           u m     ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                   �#     ����t� xa	    <�     J   J   ��     xa	J                  2         �                 � � �           u m     ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                   �#     ����t� xa	    <�     J   J   ��     xa	J                  2         �                 � � �           u m     ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                   �#     ����t� xa	    <�     J   J   ��     xa	J                  2         �                 � � �           u m     ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                   �#     ����t� xa	    <�     J   J   ��     xa	J                  2         �                 � � �           u m     ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                   �#     ����t� xa	    <�     J   J   ��     xa	J                  2         �                 � � �           u m     ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                   �#     ����t� xa	    <�     J   J   ��     xa	J                  2         �                 � � �           u m     ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                   �#     ����t� xa	    <�     J   J   ��     xa	J                  2         �                 � � �           u m     ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                   �#     ����t� xa	    <�     J   J   ��     xa	J                  2         �                 � � �           u m     ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                   �#     ����t� xa	    <�     J   J   ��     xa	J                  2         �                 � � �           u m     ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                   �#     ����t� xa	    <�     J   J   ��     xa	J                  2         �                 � � �           u m     ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                   �#     ����t� xa	    <�     J   J   ��     xa	J                  2         �                 � � �           u m     ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                   �#     ����t� xa	    <�     J   J   ��     xa	J                  2         �                 � � �           u m     ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                   �#     ����t� xa	    <�     J   J   ��     xa	J                  2         �                 � � �           u m     ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                   �#     ����t� xa	    <�     J   J   ��     xa	J                  2         �                 � � �           u m     ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                   �#     ����t� xa	    <�     J   J   ��     xa	J                  2         �                 � � �           u m     ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                   �#     ����t� xa	    <�     J   J   ��     xa	J                  2         �                 � � �           u m     ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                   �#     ����t� xa	    <�     J   J   ��     xa	J                  2         �                 � � �           u m     ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                   �#     ����t� xa	    <�     J   J   ��     xa	J                  2         �                 � � �           u m     ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                   �#     ����t� xa	    <�     J   J   ��     xa	J                  2         �                 � � �           u m     ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                               �� 	 CTitleBox                                                     �	                  $�         �  @                  ���                                                  �  @  &�     <   �  <     ��                                                        &�     |   �  |     ��    ����                                                &�     �   �  �     ��    ����                                                &�     �   �  �     ��                                                        *� h      t  4     ��                                                      h      t  4   h      t  4   [title]                                       *� �   H   �  x     ��                                                      �   H   �  x   �   H   �  x   [description]                                       *� P   �   X  �     ��                                                      P   �   X  �   P   �   X  �   [id]                                       *� �   �   �  �     ��                                                      �   �   �  �   �   �   �  �   
[designer]                                       *�      ]   1    ��        	                                                   ]   1       ]   1  Date :       �	  4  �
  �                  *� p     x  4   	 ��        
                                              p     x  4  p     x  4  [date]                                       *�       U   1    
 ��                                                            U   1         U   1   Title :       �	  4  �
  �                  *�    L   �   q     ��                                                         L   �   q      L   �   q   Description :       �	  �  �  �                  *�    �   8   �     ��                                                         �   8   �      �   8   �   ID :       �	  �  8
  J                  *�    �   �   �     ��                                                         �   �   �      �   �   �   
Designer :       �	  t  p  
                   ��������������          �     	title box     Miscellaneous      �?    9 
 ��  CParamSubBehavior    
 �  ����        ���������  ����       ���������  ����       ���������  ����       ���������  ����       ���������  ����       ���������  ����       ���������  ����       ���������  ����       ���������  ����  	     ��������        9                      �               ������   CParamSubModelType�� ����  
   ��  	 CParmDefn            title                ʃ            description                ʃ            id                ʃ            designer                ʃ            Date :                ʃ            date                ʃ            Title :                ʃ            Description :                ʃ            ID :                ʃ            
Designer :                            ����             `         �?�� 	 CGraphDoc�  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                        ���     ��   ��       ���� �        ��� 0��    2               2         �                 � � �           2       ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                         In1U2Out1Out2Out3Out4                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              1m  0                            100   100                                                           1m  0                            100   100                              1m  0                            100   100                              1m  0                            100   100                                                 
               1m  0                            100   100                            ��   CPartPackage<�T ��   CPackage@  DO14�14 pin small outline package                                                                                                                                                                                                                              ����   ������   ׃�GU ك@  DO14�14 pin small outline package                                                                                                                                                                                                                              ����   ������   ׃D�X ك@  DO14�14 pin small outline package                                                                                                                                                                                                                              ����   ������   ׃     ك�   DIP-14�14 pin dual in line package                                                                                                                                                                                                                               �     ����������������   � ��   CMiniPartPin    ����JJ     INJ�      �   ����CkCk     INCk�     �   ����KK     INK�     �   ����RR     INR�     �   ����QQ     OUTQ�     �   ����Q'Q'     OUTQ'�          ��   CPackagePin 10 RIN 
 BB.R� 1 JIN  AJ� 4 KIN  AK� 8 JIN  BB.J� 11 KIN  BB.K� 3 QOUT  AA.Q� 2 Q'OUT  AA.Q'� 13 RIN  AA.R� 5 QOUT  BB.Q� 6 Q'OUT  BB.Q'� 9 CkIN 	 BB.Clk� 12 CkIN  AA.ClkJK Flip-Flop w/clear
Flip FlopsGenericC      74107 A74107DA1               DIP1474107D74107D��  CXSpiceBehavior       jkclkresetoutnout ��   CBehPin     j����    �  j����                         ����    k����   �  k����                         ����    clk����   �  clk����                         ����     set����   �  set����                         ����    reset����   �  reset����                         ����    out����   �  out����                        ����    nout����   �  nout����                        ��74107 (XSpice)74107 (XSpice)  8               �������Digital<   Generic               ����    * time value noutQ'jJkKresetRoutQclkCk CkclkJjKkQ'noutQoutRreset                                                     � �    ����JJ     INJ�      �   ����CkCk     INCk�     �   ����KK     INK�     �   ����RR     INR�     �   ����QQ     OUTQ�     �   ����Q'Q'     OUTQ'�          ������������JK Flip-Flop w/clear
Flip FlopsGenericC      74107 A74107DA1               DIP1474107D74107D��       jkclkresetoutnout ��     j����    �  j����                         ����    k����   �  k����                         ����    clk����   �  clk����                         ����     set����   �  set����                         ����    reset����   �  reset����                         ����    out����   �  out����                        ����    nout����   �  nout����                        ��74107 (XSpice)74107 (XSpice)  8               	
Digital<   Generic               ����    * time value noutQ'jJkKresetRoutQclkCk CkclkJjKkQ'noutQoutRreset                                                     � �    ����JJ     INJ�      �   ����CkCk     INCk�     �   ����KK     INK�     �   ����RR     INR�     �   ����QQ     OUTQ�     �   ����Q'Q'     OUTQ'�       <   � 10 RIN 
 BB.R� 1 JIN  AJ� 4 KIN  AK� 8 JIN  BB.J� 11 KIN  BB.K� 3 QOUT  AA.Q� 2 Q'OUT  AA.Q'� 13 RIN  AA.R� 5 QOUT  BB.Q� 6 Q'OUT  BB.Q'� 9 CkIN 	 BB.Clk� 12 CkIN  AA.ClkJK Flip-Flop w/clear
Flip FlopsGenericC      74107 A74107DA2               DIP1474107D74107D��       jkclkresetoutnout ��     j����    �  j����                         ����    k����   �  k����                         ����    clk����   �  clk����                         ����     set����   �  set����                         ����    reset����   �  reset����                         ����    out����   �  out����                        ����    nout����   �  nout����                        ��74107 (XSpice)74107 (XSpice)  8                !"#$%&Digital<   Generic               ����    * time value noutQ'jJkKresetRoutQclkCk CkclkJjKkQ'noutQoutRreset                                                     � �    ����JJ     INJ�      �   ����CkCk     INCk�     �   ����KK     INK�     �   ����RR     INR�     �   ����QQ     OUTQ�     �   ����Q'Q'     OUTQ'�       <   JK Flip-Flop w/clear
Flip FlopsGenericC      74107 A74107DA2               DIP1474107D74107D��       jkclkresetoutnout ��     j����    �  j����                         ����    k����   �  k����                         ����    clk����   �  clk����                         ����     set����   �  set����                         ����    reset����   �  reset����                         ����    out����   �  out����                        ����    nout����   �  nout����                        ��74107 (XSpice)74107 (XSpice)  8               ./01234Digital<   Generic               ����    * time value noutQ'jJkKresetRoutQclkCk CkclkJjKkQ'noutQoutRreset                                                        �    ����AA     INA      InputInput                  �    ����AA     INA�      ClockClock               � �    ����inIn     PAS1A�      �   ����outY     PAS1Y�      '  � 1 inPAS  A1A� 2 outPAS  A1Y� 3 inPAS  B2A� 4 outPAS  B2Y� 5 inPAS  C3A� 6 outPAS  C3Y� 7  GND  COMGND� 8 outPAS  D4Y� 9 inPAS 	 D4A� 10 outPAS 
 E5Y� 11 inPAS  E5A� 12 outPAS  F6Y� 13 inPAS  F6A� 14  VCC  COMVCCdigital one-bit-wide inverterGatesGeneric=      7404 A7404DA3                                DIP147404D7404D��       inout ��     in����    �  in����                         ����    out����   �  out����                        ��7404 LS Inverter7404 LS Inverter  8               HIDigital<   Generic               ����    * time value inInoutY IninYout                        �    ����portport       ��������Output_PortOutput_Port                  �    ����portport       ��������Output_PortOutput_Port                  �    ����portport       ��������Output_PortOutput_Port                  �    ����portport       ��������Output_PortOutput_Port               � �    ����aA     IN1A�  �C  �   ����bB     IN1B�  �C  �   ����yY     OUT1Y�  �C      � 1 a   A1A� 2 b   A1B� 3 y   A1Y� 4 a   B2A� 5 b   B2B� 6 y   B2Y� 7  GND  COMGND� 8 y   C3Y� 9 a  	 C3A� 10 b  
 C3B� 11 y   D4Y� 12 a   D4A� 13 b   D4B� 14  VCC  COMVCCquad 2-input xor gatesGatesGeneric=      7486 A74LS86NA4                        DIP1474LS86N74LS86N��       aby �� �C  a����    (  a����                        ���� �C  b����   (  b����                        ���� �C  y����   (  y����                        ��74LS86 (XSpice)74LS86 (XSpice)  8               `abDigital<   Generic                       * time value yYaAbB YyAaBb                                                                       