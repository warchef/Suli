    � B2SPICE zzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzz    ��  CPart          @           @                 74107D��  CIntPin    ��  CWire      �        �       �   �  p      �   �  p              74LS08N�    �	    �   
  	 �         @           @                 74107D�    �     �       �
       �   �  p      �   �  p              74ALS11A�    
  	  25 �   �    �       24  �       24  ��  	 TModelPin    Q'����   ����Q'����                         �� �  :�0�ye>40ns��    ��������      x��    �������� �   I�����Z>25ns��    �������� �   I�����Z>25ns��    ��������      x��    �������� �   ��&�.Q>16ns��    �������� d   :�0�yE>10e-9��    �������� d   :�0�yE>10e-9��    ��������                           ����  ����:�0�yE>10e-9��d         ����  ����:�0�yE>10e-9��d   �      ��   TJKFF_general       JCkKRQQ' �     J����    ����J����                          ��      x��    ��������      x��    ��������      x��    ��������      x��    ��������      x��    ��������      x��    �������� d   :�0�yE>10e-9��    �������� d   :�0�yE>10e-9��    ��������                             ����  ����:�0�yE>10e-9��d         ����  ����:�0�yE>10e-9��d   �         �����     ��   d   :�0�yE>10e-9��    �������� d   :�0�yE>10e-9��    ���������    Ck����   ����Ck����                          ��      x��    ��������      x��    ��������      x��    ��������      x��    ��������      x��    ��������      x��    �������� d   :�0�yE>10e-9��    �������� d   :�0�yE>10e-9��    ��������                            ����  ����:�0�yE>10e-9��d         ����  ����:�0�yE>10e-9��d   �     �    �       11 �      �         @           @                 74107D�    �
      �   !   
 �       �   �  p      �   �  p              74LS08N�    �    �   %    19 $ �    %    ��   TOutPort       _   @         _   @                 Output_Port' ��  CExtPin    ��  CVertex   �  �   ��  CSegment(   - ,�?   �  �   .�*   ,�#   �  �   .�#   2 ,�   �  �   3            1     0     .�"   ,�!   @  �   5 .�!   6 ,�    @  �   7 .�    ,�   �  �   9 .�   : ,�+   �  �   ;                8                 0     /                        �   port     �  �          Q0     ��   CPin                   ��                                                           @   port�� 
 TRectangle         �   `                   ����                                                 �   `   ��  TLine     @       @      ��                                                        ��  TEllipse    8       H                  ����
[negative]               ���                       8       H      8       H   ��  
 TTextField (   ,   :   Q     ��                                                      (   ,   :   Q   (   ,   :   Q   [value]       X  d  �  �  (   ,   �   T   E�     $       <     ��                                                           $       <       $       <   [port.nbits]      <       ����            �      "Arial                    $       <   E�     ����M         ��                                                           ����M           ����M       	[refname]       @  �  �  h      �����       B   > D F G H @      Output_Port     Miscellaneous      �?      ��   TOutPortModel       port � ����port����        port����                                         0��    ��������             0��    ��������             0��    ��������             0��    ��������             0��    ��������             0��    �������� d   :�0�yE>10e-9��    �������� d   :�0�yE>10e-9��    ��������                             ����  ����:�0�yE>10e-9��d         ����  ����:�0�yE>10e-9��d   �     % J   �����     ��   d   :�0�yE>10e-9��    �������� d   :�0�yE>10e-9��    ��������Output_PortOutput_Port   �            K Digital<   Generic   Q0Q0           ����  ��    �������� ����  ��    �������� ����  ��    �������� ����  ��    �������� ����  ��    �������� ����  ��    �������� ����  ��    ��������          ����       ����  Out ��   CPartPin    ����portport       A �>      Digital Instruments Generic                                                                                                             19  K �    Q����   ����Q����                         �� �  :�0�ye>40ns��    ��������      x��    �������� �   I�����Z>25ns��    �������� �   I�����Z>25ns��    ��������      x��    �������� �   ��&�.Q>16ns��    �������� d   :�0�yE>10e-9��    �������� d   :�0�yE>10e-9��    ��������                            ����  ����:�0�yE>10e-9��d         ����  ����:�0�yE>10e-9��d   �     % �       JCkKRQQ' �     J����    ����J����                          ��      x��    ��������      x��    ��������      x��    ��������      x��    ��������      x��    ��������      x��    �������� d   :�0�yE>10e-9��    �������� d   :�0�yE>10e-9��    ��������                             ����  ����:�0�yE>10e-9��d         ����  ����:�0�yE>10e-9��d   �     ! O   �����     ��   d   :�0�yE>10e-9��    �������� d   :�0�yE>10e-9��    ���������    Ck����   ����Ck����                          ��      x��    ��������      x��    ��������      x��    ��������      x��    ��������      x��    ��������      x��    �������� d   :�0�yE>10e-9��    �������� d   :�0�yE>10e-9��    ��������                            ����  ����:�0�yE>10e-9��d         ����  ����:�0�yE>10e-9��d   �      O   �����     ��   d   :�0�yE>10e-9��    �������� d   :�0�yE>10e-9��    ���������    K����   ����K����                          ��      x��    ��������      x��    ��������      x��    ��������      x��    ��������      x��    ��������      x��    �������� d   :�0�yE>10e-9��    �������� d   :�0�yE>10e-9��    ��������                             ����  ����:�0�yE>10e-9��d         ����  ����:�0�yE>10e-9��d   �     �    �   S    14 �    S    ��   TInPort       _   @         _   @                 InputU *�    ,�   �  �   .�   Y ,�    �  `   Z .�   [ ,�   @  `   \ .�   ] ,�U   �  `   ^                                       @  �   A    �             In4     =�                    ��                                                       �   @   AC� �   8   �   H                  ����
[negative]               ���                    �   8   �   H   �   8   �   H   ?� t       �   @                   ����A                                      t       �   @   ?� t   @   �   `                   ����A                                      t   @   �   `   A� �   @   �   @     ��     	                                                  ?�         �   `                   ����                                                 �   `   A� t       t   `     
 ��                                                     ��  TPolygon                    ��                                                       ��  TPoint�   \       i��   P       i��   P       i��   D       i��   D    `  i��   P       i��   P    `yW    g�                    ��                                                       i��   $       i��   0    `  i��   0        i��   <       i��   <    �  i��   0    �  i��   0    `xW    E� �       �   8    	 ��        	                                               �       �   8   �       �   8   	[A.nbits]      <       ����            �      "Arial                �       �   8   E�    (      M     ��        
                                                 (      M      (      M   [value]       �  �  �  .     (   l   P   E� ��������+   #     ��                                                       ��������+   #   ��������+   #   	[refname]       �    "  �  ���������       ` e   d   c q   z h y { b   a f      input_general     Miscellaneous      �?      ��   TInPortModel       A �     A����    ����A����                         ��             0��    ��������             0��    ��������             0��    ��������             0��    ��������             0��    ��������             0��    �������� d   :�0�yE>10e-9��    �������� d   :�0�yE>10e-9��    ��������                            ����  ����:�0�yE>10e-9��d         ����  ����:�0�yE>10e-9��d   �     S }   �����        d   :�0�yE>10e-9��    �������� d   :�0�yE>10e-9��    ��������1 Bit Inport1 Bit Inport   �t            ~ Digital<   Generic   In4In4           ����  ��    �������� ����  ��    �������� ����  ��    �������� ����  ��    �������� ����  ��    �������� ����  ��    �������� ����  ��    ��������          ����            In L�    ����AA      INAA�?  ����Digital Instruments Generic                         `   `              `   �  �              `   �             �  `   `          �      14  R ~  14O   �����     ��   d   :�0�yE>10e-9��    �������� d   :�0�yE>10e-9��    ���������    R����   ����R����                          ��      x��    ��������      x��    ��������      x��    ��������      x��    ��������      x��    ��������      x��    �������� d   :�0�yE>10e-9��    �������� d   :�0�yE>10e-9��    ��������                            ����  ����:�0�yE>10e-9��d         ����  ����:�0�yE>10e-9��d   �     �    �   �    22 �    �    V�	       _   @         _   @                 Input� *�    ,�   @      .�C   ,�P   @  �   � .�   ,�      �   �        �         �     .�   � ,�O   �      .�   ,�@      �   �         �     � .�   � ,�G   �      � .�   ,�W   �      � .�   ,�N   `      �        �         �                        	        @  �   A      @          In1     =�                    ��                                                       �   @   AC� �   8   �   H                  ����
[negative]               ���                    �   8   �   H   �   8   �   H   ?� t       �   @                   ����A                                      t       �   @   ?� t   @   �   `                   ����A                                      t   @   �   `   A� �   @   �   @     ��                                                        ?�         �   `                   ����                                                 �   `   A� t       t   `     
 ��                                                      g�                    ��                                                       i��   \       i��   P       i��   P       i��   D       i��   D    `  i��   P       i��   P    `yW    g�                    ��                                                       i��   $       i��   0    `  i��   0        i��   <       i��   <    �  i��   0    �  i��   0    `xW    E� �       �   8    	 ��        	                                               �       �   8   �       �   8   	[A.nbits]      <       ����            �      "Arial                �       �   8   E�    (      M     ��        
                                                 (      M      (      M   [value]         �  D  N     (   l   P   E� ��������+   #     ��                                                       ��������+   #   ��������+   #   	[refname]       �  1  �  �  ���������       � �   �   � �   � � � � �   � �      input_general     Miscellaneous      �?      |�       A �     A����    ����A����                         ��             0��    ��������             0��    ��������             0��    ��������             0��    ��������             0��    ��������             0��    �������� d   :�0�yE>10e-9��    �������� d   :�0�yE>10e-9��    ��������                            ����  ����:�0�yE>10e-9��d         ����  ����:�0�yE>10e-9��d   �     � �   �����        d   :�0�yE>10e-9��    �������� d   :�0�yE>10e-9��    ��������1 Bit Inport1 Bit Inport   �t            � Digital<   Generic   In1In1           ����  ��    �������� ����  ��    �������� ����  ��    �������� ����  ��    �������� ����  ��    �������� ����  ��    �������� ����  ��    ��������  Lo�    ����            In L�    ����AA      INAAQ  ����Digital Instruments Generic                         `   `              `   �  �              `   �             �  `   `          �      22 �   �    22 �   �    22  �    R����   ����R����                          ��      x��    ��������      x��    ��������      x��    ��������      x��    ��������      x��    ��������      x��    �������� d   :�0�yE>10e-9��    �������� d   :�0�yE>10e-9��    ��������                            ����  ����:�0�yE>10e-9��d         ����  ����:�0�yE>10e-9��d   �     �    �����     ��   d   :�0�yE>10e-9��    �������� d   :�0�yE>10e-9��    ���������    R����   ����R����                          ��      x��    ��������      x��    ��������      x��    ��������      x��    ��������      x��    ��������      x��    �������� d   :�0�yE>10e-9��    �������� d   :�0�yE>10e-9��    ��������                            ����  ����:�0�yE>10e-9��d         ����  ����:�0�yE>10e-9��d   �     � �       JCkKRQQ' �     J����    ����J����                          ��      x��    ��������      x��    ��������      x��    ��������      x��    ��������      x��    ��������      x��    �������� d   :�0�yE>10e-9��    �������� d   :�0�yE>10e-9��    ��������                             ����  ����:�0�yE>10e-9��d         ����  ����:�0�yE>10e-9��d   �      �   �����     ��   d   :�0�yE>10e-9��    �������� d   :�0�yE>10e-9��    ���������    Ck����   ����Ck����                          ��      x��    ��������      x��    ��������      x��    ��������      x��    ��������      x��    ��������      x��    �������� d   :�0�yE>10e-9��    �������� d   :�0�yE>10e-9��    ��������                            ����  ����:�0�yE>10e-9��d         ����  ����:�0�yE>10e-9��d   �      �   �����     ��   d   :�0�yE>10e-9��    �������� d   :�0�yE>10e-9��    ���������    K����   ����K����                          ��      x��    ��������      x��    ��������      x��    ��������      x��    ��������      x��    ��������      x��    �������� d   :�0�yE>10e-9��    �������� d   :�0�yE>10e-9��    ��������                             ����  ����:�0�yE>10e-9��d         ����  ����:�0�yE>10e-9��d   �     �    �   �    9 �    �    V�       _   @         _   @                 Input� *�    ,�   `      .�H   � ,�   �      �                       @  �   A       @          In2     =�                    ��                                                       �   @   AC� �   8   �   H                  ����
[negative]               ���                    �   8   �   H   �   8   �   H   ?� t       �   @                   ����A                                      t       �   @   ?� t   @   �   `                   ����A                                      t   @   �   `   A� �   @   �   @     ��    ����                                                ?�         �   `                   ����                                                 �   `   A� t       t   `     
 ��                                                      g�                    ��                                                       i��   \       i��   P       i��   P       i��   D       i��   D    `  i��   P       i��   P    `yW    g�                    ��                                                       i��   $       i��   0    `  i��   0        i��   <       i��   <    �  i��   0    �  i��   0    `xW    E� �       �   8    	 ��        	                                               �       �   8   �       �   8   	[A.nbits]      <       ����            �      "Arial                �       �   8   E�    (      M     ��        
                                                 (      M      (      M   [value]       ,  �  d  N     (   l   P   E� ��������+   #     ��                                                       ��������+   #   ��������+   #   	[refname]         1  �  �  ���������       � �   �   � �   � � � � �   � �      input_general     Miscellaneous      �?      |�       A �     A����    ����A����                         ��             0��    ��������             0��    ��������             0��    ��������             0��    ��������             0��    ��������             0��    �������� d   :�0�yE>10e-9��    �������� d   :�0�yE>10e-9��    ��������                            ����  ����:�0�yE>10e-9��d         ����  ����:�0�yE>10e-9��d   �     � �   �����        d   :�0�yE>10e-9��    �������� d   :�0�yE>10e-9��    ��������1 Bit Inport1 Bit Inport   �t            � Digital<   Generic   In2In2           ����  ��    �������� ����  ��    �������� ����  ��    �������� ����  ��    �������� ����  ��    �������� ����  ��    �������� ����  ��    ��������  4�    ����            In L�    ����AA      INAA�?  ����Digital Instruments Generic                         `   `              `   �  �              `   �             �  `   `          �      9  � �  9�   �����     ��   d   :�0�yE>10e-9��    �������� d   :�0�yE>10e-9��    ��������� �    Q����   ����Q����                         �� �  :�0�ye>40ns��    ��������      x��    �������� �   I�����Z>25ns��    �������� �   I�����Z>25ns��    ��������      x��    �������� �   ��&�.Q>16ns��    �������� d   :�0�yE>10e-9��    �������� d   :�0�yE>10e-9��    ��������                            ����  ����:�0�yE>10e-9��d         ����  ����:�0�yE>10e-9��d   �     �    �   �    13 �    �    (�       _   @         _   @                 Output_Port� *�    ,�      �   .�I   � ,�V      �   � .�G   � ,�T   �  �   � .�F   � ,�H   �  @   � .�B   ,�      @   .�D   ,�D   �  @   �     �     �        �                                            �   port                   Q2     =�                   ��                                                           @   port?�         �   `                   ����                                                 �   `   A�     @       @      ��                                                        C�    8       H                  ����
[negative]               ���                       8       H      8       H   E� (   ,   :   Q     ��                                                      (   ,   :   Q   (   ,   :   Q   [value]       x  �  �    (   ,   �   T   E�     $       <     ��                                                           $       <       $       <   [port.nbits]      <       ����            �      "Arial                    $       <   E�     ����M         ��                                                           ����M           ����M       	[refname]       `  �  �  �      �����       �   � � � � � �      Output_Port     Miscellaneous      �?      I�       port � ����port����        port����                                         0��    ��������             0��    ��������             0��    ��������             0��    ��������             0��    ��������             0��    �������� d   :�0�yE>10e-9��    �������� d   :�0�yE>10e-9��    ��������                             ����  ����:�0�yE>10e-9��d         ����  ����:�0�yE>10e-9��d   �     � �   �����     ��   d   :�0�yE>10e-9��    �������� d   :�0�yE>10e-9��    ��������Output_PortOutput_Port                 � Digital<   Generic   Q2Q2           ����  ��    �������� ����  ��    �������� ����  ��    �������� ����  ��    �������� ����  ��    �������� ����  ��    �������� ����  ��    ��������          ����       ����  Out L�    ����portport       A ����    Digital Instruments Generic                                                                                                             13  � �  13�   �����         d   :�0�yE>10e-9��    �������� d   :�0�yE>10e-9��    ���������    Q'����   ����Q'����                         �� �  :�0�ye>40ns��    ��������      x��    �������� �   I�����Z>25ns��    �������� �   I�����Z>25ns��    ��������      x��    �������� �   ��&�.Q>16ns��    �������� d   :�0�yE>10e-9��    �������� d   :�0�yE>10e-9��    ��������                           ����  ����:�0�yE>10e-9��d         ����  ����:�0�yE>10e-9��d   �     
 �   �����        d   :�0�yE>10e-9��    �������� d   :�0�yE>10e-9��    ��������107 JK FF w/clear107 JK FF w/clear   �t            � � � � � � Digital<   Generic   A1A1           ���� x��    �������� ���� x��    �������� �'	 hUMu?60u��    �������� ʑ�b2U0*�c�-2.4m��    �������� ���-C��6:�-.4m��    ��������  h�	����Mb�?16m��    ��������  ��{�G�z�?10m��    ��������          ����Standard TTL                 0��    �������� ����    �sA20meg��    �������� 6  ��创�`>31n��    ��������             0��    ��������  �����     ��   d   :�0�yE>10e-9��    �������� d   :�0�yE>10e-9��    ��������� �  22O   �����     ��   d   :�0�yE>10e-9��    �������� d   :�0�yE>10e-9��    ��������N �    Q'����   ����Q'����                         �� �  :�0�ye>40ns��    ��������      x��    �������� �   I�����Z>25ns��    �������� �   I�����Z>25ns��    ��������      x��    �������� �   ��&�.Q>16ns��    �������� d   :�0�yE>10e-9��    �������� d   :�0�yE>10e-9��    ��������                           ����  ����:�0�yE>10e-9��d         ����  ����:�0�yE>10e-9��d   �     �    �   �    26 �   �    26  � �    C����   ����C����                          ��      x��    ��������      x��    ��������      x��    ��������      x��    ��������      x��    ��������      x��    �������� d   :�0�yE>10e-9��    �������� d   :�0�yE>10e-9��    ��������                             ����  ����:�0�yE>10e-9��d         ����  ����:�0�yE>10e-9��d   �     � ��   TAnd       ABCY �     A����    ����A����                          ��      x��    ��������      x��    ��������      x��    ��������      x��    ��������      x��    ��������      x��    �������� d   :�0�yE>10e-9��    �������� d   :�0�yE>10e-9��    ��������                             ����  ����:�0�yE>10e-9��d         ����  ����:�0�yE>10e-9��d   �     
   �����     ��   d   :�0�yE>10e-9��    �������� d   :�0�yE>10e-9��    ���������    B����   ����B����                          ��      x��    ��������      x��    ��������      x��    ��������      x��    ��������      x��    ��������      x��    �������� d   :�0�yE>10e-9��    �������� d   :�0�yE>10e-9��    ��������                             ����  ����:�0�yE>10e-9��d         ����  ����:�0�yE>10e-9��d   �        �����     ��   d   :�0�yE>10e-9��    �������� d   :�0�yE>10e-9��    ��������� �    Y����   ����Y����                         �� d   :�0�yE>10ns��    ��������    ��&�.!>2ns��    ��������      x��    �������� �   �?Y��K>13ns��    ��������    ��&�.!>2ns��    ��������      x��    �������� d   :�0�yE>10e-9��    �������� d   :�0�yE>10e-9��    ��������                            ����  ����:�0�yE>10e-9��d         ����  ����:�0�yE>10e-9��d   �        �����        d   :�0�yE>10e-9��    �������� d   :�0�yE>10e-9��    ��������11A/3 ALS 3-input And11A/3 ALS 3-input And  D �t            � Digital<   Motorola   U3U3           ���� x��    �������� ���� x��    �������� @ �h㈵��>20u��    �������� ����-C��6�-.1m��    �������� ���-C��6:�-.4m��    ��������  ������Mb�?8m��    �������� @]� ��_�LU?1.3m��    ��������         ����ALS      �����     ��   d   :�0�yE>10e-9��    �������� d   :�0�yE>10e-9��    �������� 26O   �����        d   :�0�yE>10e-9��    �������� d   :�0�yE>10e-9��    ��������107 JK FF w/clear107 JK FF w/clear   �            P Q R � N � Digital<   Generic   A3A3           ���� x��    �������� ���� x��    �������� �'	 hUMu?60u��    �������� ʑ�b2U0*�c�-2.4m��    �������� ���-C��6:�-.4m��    ��������  h�	����Mb�?16m��    ��������  ��{�G�z�?10m��    ��������          ����Standard TTL                 0��    �������� ����    �sA20meg��    �������� 6  ��创�`>31n��    ��������             0��    ��������  �����         d   :�0�yE>10e-9��    �������� d   :�0�yE>10e-9��    ��������� ;  A����        A����                          ��      x��    ��������      x��    ��������      x��    ��������      x��    ��������      x��    ��������      x��    �������� d   :�0�yE>10e-9��    �������� d   :�0�yE>10e-9��    ��������                             ����  ����:�0�yE>10e-9��d         ����  ����:�0�yE>10e-9��d   �     %  �       ABY � <  B����       B����                          ��      x��    ��������      x��    ��������      x��    ��������      x��    ��������      x��    ��������      x��    �������� d   :�0�yE>10e-9��    �������� d   :�0�yE>10e-9��    ��������                             ����  ����:�0�yE>10e-9��d         ����  ����:�0�yE>10e-9��d   �        �����     ��   d   :�0�yE>10e-9��    �������� d   :�0�yE>10e-9��    ��������� =  Y����       Y����                         �� �   :�0�yU>20ns��    ��������      x��    �������� d   :�0�yE>10ns��    �������� �   ,i�)+P>15ns��    ��������      x��    �������� P   ��&�.A>8ns��    �������� d   :�0�yE>10e-9��    �������� d   :�0�yE>10e-9��    ��������                            ����  ����:�0�yE>10e-9��d         ����  ����:�0�yE>10e-9��d   �     !   �����         d   :�0�yE>10e-9��    �������� d   :�0�yE>10e-9��    ��������08/4 LS 2-Inp. And08/4 LS 2-Inp. And  A �t            Digital<   Analog Devices   A5A5           ���� x��    �������� ���� x��    �������� @ �h㈵��>20u��    �������� ���-C��6:�-.4m��    �������� ���-C��6:�-.4m��    ��������  ������Mb�?8m��    �������� ��`�Q�k?3.4m��    ��������          ����LS      �����     ��   d   :�0�yE>10e-9��    �������� d   :�0�yE>10e-9��    �������� 19  # 19 �       # 1 " *�    ,�-   �  @   .�   ,�   �  �   .�   ,�   @  �   .�   ,�   �  �    
        
            
        
         �  �  y    *�   <           a   *�   ,�*   �  �   .�$   ,�&      �   .�&   ,�(          .�)   ,�E   �
      .�5   ,�;   �
  @   .�4   ,�      @   .�3   ,�:   `  @                                                                                �  b    �  �          A5     =�                   ��                                                       �   �   y=�                    ��                                                          `   a=�                   ��                                                          �   bA�     P       �    
 ��    ��W                                                A�     �       �    	 ��    x��                                                A�     `       `     ��    ����                                                A� �   �   �   �     ��                                                       A�     �   D   �     ��    �U �                                                ��   TArc    P   �   �                                                                  P   �   �      P   �   �   �   �   D   P           A�     P   D   P     ��     	  	                                                )�    0   �   �               
                                                   0   �   �      0   �   �   D   �   �   �           E�     �����        ��                                                           �����          �����      	[devname]        ����������������    �����      E�        b   D     ��                                                              b   D          b   D   	[refname]            �  �         �   @    "#  ,  +!*  (  .'-  &  %  $     AND 2    
AND 2 IEEEMiscellaneous      �?    A    A L�    ����aA      INA1A�?      L�   ����bB      INA1B�?     L�   ����yY      OUTA1Y�?     L�    ����aA      INB1A�?      L�   ����bB      INB1B����   L�   ����yY      OUTB1Y�?     L�    ����aA      INC1A�?      L�   ����bB      INC1B�?     L�   ����yY      OUTC1Y       L�    ����aA      IND1A�?      L�   ����bB      IND1B�?     L�   ����yY      OUTD1Y       GatesXSpice 2input AND gateGenericDIP-14             15  P 
 15  
  15  T � & � *�           �  J�  *�   ,�
   @      .�   ,�   �      .�   ?,�"   �  `	   .�	   ,�2   �  `	   .�   ,�%   �  �   D.�
   E,�      �   F                C    B.�   ,�K      `	   .�'   ,�<      �   J.�%   ,�9   �  �   L.�   ,�8   �  �   N.�   O,�   �  �   P.�   Q,�6   @  �   R                       M        K        I    H        C        A    @        >    =    .�   =,�   �      T                     �  Ck�  *�   ]       @  K�  *�   �         R�  *�   4   @  �  Q�  *�   ,�   �  `   .�8   Z,�I   �  `   [.�7   ,�F   �  `    ].�6   ,�)          _   
    ^        \                     @  @  Q'�   @             A3     =�                    ��                                                           �   J=�                   ��                                                          �   Ck=�                   ��                                                          �   K=�                   ��                                                      `      R=�                   ��                                                      �   �   Q=�                   ��                                                      �   �   Q'?�     `   �   �                  ����                                             `   �   �   A�     �       �     ��                                                        A�     �       �     ��                                                        A�     �       �    	 ��        	                                                A� `   �   `       
 ��    ����
                                                A� �   �   �   �     ��    ����                                                A� �   �   �   �     ��    ����                                                A� �   x   �   �     ��    ����                                                A� �   x   �   x     ��    ����                                                C� X   �   h   �                  �                                           X   �   h   �   X   �   h   �   A� �   �   �   �     ��    ����                                                A� �   �   �   �     ��    ����                                                C� �   �   �   �                  �                                           �   �   �   �   �   �   �   �   E�     0   b   X     ��                                                           0   b   X       0   b   X   	[refname]       �  �  h  P      0   �   T   E� (   p   0   �     ��                                                      (   p   0   �   (   p   0   �   j       �  p  �    (   p   p   �   E� (   �   P   �     ��                                                      (   �   P   �   (   �   P   �   clk       �  �  0  f  (   �   p   �   E� (   �   8   �     ��                                                      (   �   8   �   (   �   8   �   k       �  0  �  �  (   �   p   �   E�        �   0     ��                                                              �   0          �   0   	[devname]        ����������������       �   0    abcdefghijklmuvw      o  qrxnst  p     74107 JK FF w/clear    74107 JK FF w/clear IEEEMiscellaneous      �?      O   A L�    ����JJ      INAJ�>  ����L�   ����CkCk      INACk�>  ����L�   ����KK      INAK�>  ����L�   ����RR      INAR�>  ����L�   ����QQ      OUTAQ�>  ����L�   ����Q'Q'      OUTAQ'��������L�    ����JJ      INBJ�>  ����L�   ����CkCk      INBCk�>  ����L�   ����KK      INBK�>  ����L�   ����RR      INBR�>  ����L�   ����QQ      OUTBQ�>  ����L�   ����Q'Q'      OUTBQ'�>  ����
Flip FlopsJK Flip-Flop w/clearGenericDO14              11 �        ��   TClock       �   �  �      �   �  �              Clock�*�    I   �     A�   `  @          U1     =�                   ��                                                       �   `   A?�     @   �   �                  ����                                             @   �   �   A� �   `   �   `     ��    �X                                                A� `   @   `   �     ��    8�W                                                A� p   h   x   h     ��    ��W                                                A� x   T   x   h     ��    X                                                A� x   T   �   T     ��    ��W                                                A� �   T   �   h     ��    �W                                                A� �   h   �   h     ��     X                                                A� �   P   �   p      ��    8�W	                                                E�    P   Z   u    
 ��        
                                                  P   Z   u      P   Z   u   [period]       �  0	  p  �	     P   P   t   E� �   `   �   �    	 ��                                                      �   `   �   �   �   `   �   �   ns       @  `	  �  �	  �   `   �   x   E�     �����        ��                                                           �����          �����      	[devname]        ����������������    �����      E�        *   @     ��                                                              *   @          *   @   	[refname]       `  �  �  (	         �   <    �  �  �  �  ��  ����  �  �  �    �     Clock     Miscellaneous      �?      ��   TClockModel     ��  CValue �  I�����z>100n      ���������� �  I�����j>50n     �������� A �     A����    ����A����                          ��      x��    ��������      x��    ��������      x��    ��������      x��    ��������      x��    ��������      x��    �������� d   :�0�yE>10e-9��    �������� d   :�0�yE>10e-9��    ��������                             ����  ����:�0�yE>10e-9��d         ����  ����:�0�yE>10e-9��d   �      �  �����         d   :�0�yE>10e-9��    �������� d   :�0�yE>10e-9��    ��������ClockClock              �Digital InstrumentsO   Generic   U1U1           ����  ��    �������� ����  ��    �������� ����  ��    �������� ����  ��    �������� ����  ��    �������� ����  ��    �������� ����  ��    ��������  al      ����Generic             U L�    ����AA      INAA�  ����Digital InstrumentsDigital Clock inputGeneric                                                                              �'                                   11 �       11   � Q � 11   �����     ��   d   :�0�yE>10e-9��    �������� d   :�0�yE>10e-9��    ���������    K����   ����K����                          ��      x��    ��������      x��    ��������      x��    ��������      x��    ��������      x��    ��������      x��    �������� d   :�0�yE>10e-9��    �������� d   :�0�yE>10e-9��    ��������                             ����  ����:�0�yE>10e-9��d         ����  ����:�0�yE>10e-9��d   �     �    �   �   3 �    �   V�       _   @         _   @                 Input�*�    ,�   @      .�   �,�   @      �.�   �,�	          �.�   �,�   `      �                                       @  �   A     	  `          In3     =�                    ��                                                       �   @   AC� �   8   �   H                  ����
[negative]               ���                    �   8   �   H   �   8   �   H   ?� t       �   @                   ����A                                      t       �   @   ?� t   @   �   `                   ����A                                      t   @   �   `   A� �   @   �   @     ��                                                        ?�         �   `                   ����                                                 �   `   A� t       t   `     
 ��                                                      g�                    ��                                                       i��   \       i��   P       i��   P       i��   D       i��   D    `  i��   P       i��   P    `yW    g�                    ��                                                       i��   $       i��   0    `  i��   0        i��   <       i��   <    �  i��   0    �  i��   0    `xW    E� �       �   8    	 ��        	                                               �       �   8   �       �   8   	[A.nbits]      <       ����            �      "Arial                �       �   8   E�    (      M     ��        
                                                 (      M      (      M   [value]       	  �  D	  n     (   l   P   E� ��������+   #     ��                                                       ��������+   #   ��������+   #   	[refname]       �  Q  �	  �  ���������       ��  �  ��  �����  ��     input_general     Miscellaneous      �?      |�       A �     A����    ����A����                         ��             0��    ��������             0��    ��������             0��    ��������             0��    ��������             0��    ��������             0��    �������� d   :�0�yE>10e-9��    �������� d   :�0�yE>10e-9��    ��������                            ����  ����:�0�yE>10e-9��d         ����  ����:�0�yE>10e-9��d   �     ��  �����        d   :�0�yE>10e-9��    �������� d   :�0�yE>10e-9��    ��������1 Bit Inport1 Bit Inport   �t            �Digital<   Generic   In3In3           ����  ��    �������� ����  ��    �������� ����  ��    �������� ����  ��    �������� ����  ��    �������� ����  ��    �������� ����  ��    ��������  al      ����            In L�    ����AA      INAA��������Digital Instruments Generic               ���        `   `              `   �  �              `   �             �  `   `          �      3  �� 3   �����     ��   d   :�0�yE>10e-9��    �������� d   :�0�yE>10e-9��    ��������� �    Q����   ����Q����                         �� �  :�0�ye>40ns��    ��������      x��    �������� �   I�����Z>25ns��    �������� �   I�����Z>25ns��    ��������      x��    �������� �   ��&�.Q>16ns��    �������� d   :�0�yE>10e-9��    �������� d   :�0�yE>10e-9��    ��������                            ����  ����:�0�yE>10e-9��d         ����  ����:�0�yE>10e-9��d   �     �    �   �   5 �    �   (�       _   @         _   @                 Output_Port�*�    ,�   �  `   .�>   �,�C   �  �   �.�=   �,�B   �  �   �.�<   �,�A   �  @   �.�.   ,�   @  @   �        �                                           �   port     �  �          Q1     =�                   ��                                                           @   port?�         �   `                   ����                                                 �   `   A�     @       @      ��                                                        C�    8       H                  ����
[negative]               ���                       8       H      8       H   E� (   ,   :   Q     ��                                                      (   ,   :   Q   (   ,   :   Q   [value]       �  $  0  �  (   ,   �   T   E�     $       <     ��                                                           $       <       $       <   [port.nbits]      <       ����            �      "Arial                    $       <   E�     ����M         ��                                                           ����M           ����M       	[refname]       �  �  h  (      �����       �  ������     Output_Port     Miscellaneous      �?      I�       port � ����port����        port����                                         0��    ��������             0��    ��������             0��    ��������             0��    ��������             0��    ��������             0��    �������� d   :�0�yE>10e-9��    �������� d   :�0�yE>10e-9��    ��������                             ����  ����:�0�yE>10e-9��d         ����  ����:�0�yE>10e-9��d   �     ��  �����     ��   d   :�0�yE>10e-9��    �������� d   :�0�yE>10e-9��    ��������Output_PortOutput_Port   �            �Digital<   Generic   Q1Q1           ����  ��    �������� ����  ��    �������� ����  ��    �������� ����  ��    �������� ����  ��    �������� ����  ��    �������� ����  ��    ��������          ����       ����  Out L�    ����portport       A X]      Digital Instruments Generic                                                                                                             5  �� 5   �����         d   :�0�yE>10e-9��    �������� d   :�0�yE>10e-9��    �������� 107 JK FF w/clear107 JK FF w/clear   �              �� � Digital<   Generic   A2A2           ���� x��    �������� ���� x��    �������� �'	 hUMu?60u��    �������� ʑ�b2U0*�c�-2.4m��    �������� ���-C��6:�-.4m��    ��������  h�	����Mb�?16m��    ��������  ��{�G�z�?10m��    ��������          ����Standard TTL                 0��    �������� ����    �sA20meg��    �������� 6  ��创�`>31n��    ��������             0��    ��������  �����        d   :�0�yE>10e-9��    �������� d   :�0�yE>10e-9��    ��������� <  B����       B����                          ��      x��    ��������      x��    ��������      x��    ��������      x��    ��������      x��    ��������      x��    �������� d   :�0�yE>10e-9��    �������� d   :�0�yE>10e-9��    ��������                             ����  ����:�0�yE>10e-9��d         ����  ����:�0�yE>10e-9��d   �       �       ABY � ;  A����        A����                          ��      x��    ��������      x��    ��������      x��    ��������      x��    ��������      x��    ��������      x��    �������� d   :�0�yE>10e-9��    �������� d   :�0�yE>10e-9��    ��������                             ����  ����:�0�yE>10e-9��d         ����  ����:�0�yE>10e-9��d   �     
 �  �����     ��   d   :�0�yE>10e-9��    �������� d   :�0�yE>10e-9��    ���������� =  Y����       Y����                         �� �   :�0�yU>20ns��    ��������      x��    �������� d   :�0�yE>10ns��    �������� �   ,i�)+P>15ns��    ��������      x��    �������� P   ��&�.A>8ns��    �������� d   :�0�yE>10e-9��    �������� d   :�0�yE>10e-9��    ��������                            ����  ����:�0�yE>10e-9��d         ����  ����:�0�yE>10e-9��d   �      �  �����        d   :�0�yE>10e-9��    �������� d   :�0�yE>10e-9��    ��������08/4 LS 2-Inp. And08/4 LS 2-Inp. And  A \            ���Digital<   Analog Devices   A4A4           ���� x��    �������� ���� x��    �������� @ �h㈵��>20u��    �������� ���-C��6:�-.4m��    �������� ���-C��6:�-.4m��    ��������  ������Mb�?8m��    �������� ��`�Q�k?3.4m��    ��������         ����LS      �����     ��   d   :�0�yE>10e-9��    �������� d   :�0�yE>10e-9��    �������� 24   24 �  *�    ,�'   @  �   .�   ,�5   �  �   �.�   �,�4   �  @   �.�   �,�   �  @   �.�   �,�3   @  @   �                                �       
           �  yC  *�   ,�,      �   .�:   ,�J   �  �   �    �    .�9   �,�M      �   .�;   �,�Q          �.�/   �,�0          �.�?   ,�$   @      �        �    .�-   �,�/      �   �.�,   ,�.    	  �   �.�+   ,�=    	  �           �        �                            �           
      �  �  bD  *�   ,�L      �   .�@   ,�R   �  �   .�A   ,�S   �      .�E   ,�           	          .�2   ,�7   �  �   
.�1   ,�>    	  �   .�0   ,�1   `	  �    	        	           	        	        	        	  
       �  �  aE  *�   `  �     cF   @             U3     =�                    ��                                                           �   y=�                   ��                                                      �   �   b=�                   ��                                                      �   �   a=�                   ��                                                      �   `   cA� �   �   �   �     ��     ~�                                                )� ����p   d   �                                                                  P   �   �      P   �   �   \   P      �           A� �   �   \   �    
 ��    h                                                  )� �����   d      	                                                              0   �   �      0   �   �      �   \   �           A� �   P   \   P     ��    ��                                                A�     �       �     ��    {  	                                                A� �   �   �   �     ��    (��
                                                A� �   `   �   `     ��       �                                                A� �   �   �   P     ��    ��                                                E�         *   H     ��                                                               *   H           *   H   	[refname]       @  `   �             �   D   E�     �����         ��                                                           �����           �����       	[devname]        ����������������    �����                           AND 3    
AND 3 IEEEMiscellaneous      �?    D    U L�    ����aA      INAaz	  ����L�   ����bB      INAb{	  ����L�   ����cC      INAc|	  ����L�   ����yY      OUTAy}	  ����Gatestriple 3-input AND gatesGeneric               23  �  23    23 �� � �  *�    �       �  J�  *�   Q      �  Ck�  *�   �       @  K�  *�   �         R�  *�   �   @  �  Q�  *�   	  @  @  Q'�   �  �          A1     =�                    ��                                                           �   J=�                   ��                                                          �   Ck=�                   ��                                                          �   K=�                   ��                                                      `      R=�                   ��                                                      �   �   Q=�                   ��                                                      �   �   Q'?�     `   �   �                  ����                                             `   �   �   A�     �       �     ��                                                        A�     �       �     ��                                                        A�     �       �    	 ��        	                                                A� `   �   `       
 ��        
                                                A� �   �   �   �     ��                                                        A� �   �   �   �     ��    ����                                                A� �   x   �   �     ��    ����                                                A� �   x   �   x     ��                                                        C� X   �   h   �                  �                                           X   �   h   �   X   �   h   �   A� �   �   �   �     ��                                                        A� �   �   �   �     ��                                                        C� �   �   �   �                  �                                           �   �   �   �   �   �   �   �   E�     0   b   X     ��                                                           0   b   X       0   b   X   	[refname]       @  P    �      0   �   T   E� (   p   0   �     ��                                                      (   p   0   �   (   p   0   �   j       X    p  �  (   p   p   �   E� (   �   P   �     ��                                                      (   �   P   �   (   �   P   �   clk       X  p  �    (   �   p   �   E� (   �   8   �     ��                                                      (   �   8   �   (   �   8   �   k       X  �  �  f  (   �   p   �   E�        �   0     ��                                                              �   0          �   0   	[devname]        ����������������       �   0    *+,-./0123456>?@      8  :;A7<=  90     74107 JK FF w/clear    74107 JK FF w/clear IEEEMiscellaneous      �?      �   A L�    ����JJ      INAJyE>����L�   ����CkCk      INACkE>1����L�   ����KK      INAK    ����L�   ����RR      INAR�<�����L�   ����QQ      OUTAQ   �����L�   ����Q'Q'      OUTAQ'�>  ����L�    ����JJ      INBJ��������L�   ����CkCk      INBCk�>  ����L�   ����KK      INBK�>  ����L�   ����RR      INBR�>  ����L�   ����QQ      OUTBQ�?  ����L�   ����Q'Q'      OUTBQ'�?  ����
Flip FlopsJK Flip-Flop w/clearGenericDO14              25  	  � �	 25 	  25   *�      �  �  y    *�             a   *�         �  b     	  �          A4     =�                   ��                                                       �   �   y=�                    ��                                                          `   a=�                   ��                                                          �   bA�     P       �    
 ��    ` �                                                A�     �       �    	 ��    &                                                   A�     `       `     ��    �                                                  A� �   �   �   �     ��    � �                                                A�     �   D   �     ��    ����                                                )�    P   �   �                                                                  P   �   �      P   �   �   �   �   D   P           A�     P   D   P     ��       	                                                )�    0   �   �               
                                                   0   �   �      0   �   �   D   �   �   �           E�     �����        ��                                                           �����          �����      	[devname]        ����������������    �����      E�        b   D     ��                                                              b   D          b   D   	[refname]       `	  �  (
  �         �   @    RS  [  ZQY  X  ]W\  V  U  T     AND 2    
AND 2 IEEEMiscellaneous      �?    A  �  A L�    ����aA      INA1A�>      L�   ����bB      INA1B�?     L�   ����yY      OUTA1Y�>     L�    ����aA      INB1A�>      L�   ����bB      INB1B      L�   ����yY      OUTB1Y      L�    ����aA      INC1A l     L�   ����bB      INC1B��(A   L�   ����yY      OUTC1Y      L�    ����aA      IND1A       L�   ����bB      IND1B@     L�   ����yY      OUTD1Y@     GatesXSpice 2input AND gateGenericDIP-14              1 	  �  1  �� 1  �� � *�           �  J�  *�   G      �  Ck�  *�   �      @  K�  *�   �         R�  *�   �  @  �  Q�  *�   �  @  @  Q'�      �          A2     =�                    ��                                                           �   J=�                   ��                                                          �   Ck=�                   ��                                                          �   K=�                   ��                                                      `      R=�                   ��                                                      �   �   Q=�                   ��                                                      �   �   Q'?�     `   �   �                  ����                                             `   �   �   A�     �       �     ��                                                        A�     �       �     ��                                                        A�     �       �    	 ��        	                                                A� `   �   `       
 ��    ���
                                                A� �   �   �   �     ��                                                        A� �   �   �   �     ��                                                        A� �   x   �   �     ��                                                        A� �   x   �   x     ��                                                        C� X   �   h   �                  �                                           X   �   h   �   X   �   h   �   A� �   �   �   �     ��    ���                                                A� �   �   �   �     ��                                                        C� �   �   �   �                  �                                           �   �   �   �   �   �   �   �   E�     0   b   X     ��                                                           0   b   X       0   b   X   	[refname]       `  P  (  �      0   �   T   E� (   p   0   �     ��                                                      (   p   0   �   (   p   0   �   j       x    �  �  (   p   p   �   E� (   �   P   �     ��                                                      (   �   P   �   (   �   P   �   clk       x  p  �    (   �   p   �   E� (   �   8   �     ��                                                      (   �   8   �   (   �   8   �   k       x  �  �  f  (   �   p   �   E�        �   0     ��                                                              �   0          �   0   	[devname]        ����������������       �   0    pqrstuvwxyz{|���      ~  ���}��  �     74107 JK FF w/clear    74107 JK FF w/clear IEEEMiscellaneous      �?         A L�    ����JJ      INAJ    ����L�   ����CkCk      INACk   ����L�   ����KK      INAK 5����L�   ����RR      INAR   ����L�   ����QQ      OUTAQ  x����L�   ����Q'Q'      OUTAQ'0e-9����L�    ����JJ      INBJ10e-����L�   ����CkCk      INBCk J�����L�   ����KK      INBK   ����L�   ����RR      INBR d ����L�   ����QQ      OUTBQ �������L�   ����Q'Q'      OUTBQ'yE>����
Flip FlopsJK Flip-Flop w/clearGenericDO14                �� �) � �  # �W      �� �  � � 
 ! S % � J I J   � � � � T.�   ,�            �    ,�   �       �        >@BFD� H� ���^ \ �Z RP��N�; 9 7 5 3 LJ/ 1  ����
_][�������� � � � � � � X X X [ Y ����	� �=�UG] �Z� � �� Q� �4 - : ?� 8 6 A2 �E�`< ����C���SOM K0 � ���� ^� � \�I�� � � �� _ � �              
 ��@ ����        ����������             0     ���������� ����      @5     ����������  ʚ;�������?.1     ����������@ ����       ���������� ����       ���������� ����       ���������� ����       ���������� ���� true
     ���������� ����  false     ��������               
                  �� ����        ���������� ����       ����������  ����       ����������@ ����       ����������@ ����       ��������               
                  �� ����        ���������� ����       ����������@ ����       ����������  ����       ���������� ����       ���������� ����       ���������� ����       ���������� ����       ���������� ����       ���������� ����       ���������� ����       ��������               
                 �� ����dec     ���������� ����     @�@1k     ���������� ����    ��.A1meg     ���������� ����       20     ���������� ���� true     ���������� ���� true     ���������� ���� true	     ���������� ����  false
     ��������               
                 ��  ����        ����������  ����       ����������  ����       ���������� ����dec     ���������� ����       ���������� ����       ���������� ����  	     ���������� ����  
     ��������               
                  	 �� ����        ���������� ����       ���������� ����       ���������� ����       ���������� ����       ���������� ����       ���������� ����       ���������� ����       ���������� ����       ��������               
                 �� ����        ���������� ����       ���������� ����       ���������� ����dec     ���������� ����       ��������               
                     ��             0      ���������� ��� ����MbP?1m     ���������� �� �h㈵��>10u     ���������� '  ���ư>1u     ���������� ���� true     ���������� ����  false     ���������� ���� true     ���������� ����  false     ��������               
                 �� ����     @�@1K      ����������  ����       ����������  ����       ����������  ����       ��������               
         ��              ��  ����        ��������              
                  ��  ����        ��������              
                                  
                 ��@ ����        ����������@ ����       ���������� ����       ���������� ����       ���������� ����       ���������� ����       ���������� ����       ���������� ����       ���������� ����       ���������� ���� true	     ���������� ����  false
     ���������� ���� true     ���������� ����  false     ��������               
                 �� ����       5      ���������� ����       5     ���������� ����       5     ���������� ����       5     ���������� ����       ���������� ����  	     ���������� ����  
     ���������� ����       ���������� ����       ���������� ����       ���������� ���� true     ����������@ ����       ����������@ ����       ���������� ����       ���������� ����       ���������� ����       ���������� ����dec     ���������� ����       ���������� ����       ���������� ����       ���������� ���� true     ���������� ���� true     ���������� ���� true     ���������� ����  false     ���������� ���� true     ���������� ����  false      ���������� ���� true!     ���������� ����  false"     ��������               
                        �� ����       5      ���������� ����       5     ���������� ����       5     ���������� ����       5     ���������� ����       ���������� ����  	     ���������� ����  
     ���������� ����       ���������� ����       ���������� ����       ���������� ���� true     ����������@ ����       ����������@ ����       ���������� ����       ���������� ����       ���������� ����       ���������� ����dec     ���������� ����       ���������� ����       ���������� ����       ���������� ���� true     ���������� ���� true     ���������� ���� true     ���������� ����  false     ���������� ���� true     ���������� ����  false      ���������� ���� true!     ���������� ����  false"     ��������               
                 �� ����       5      ���������� ����       5     ���������� ����       5     ���������� ����       5     ���������� ����       ���������� ����  	     ���������� ����  
     ���������� ����       ���������� ����       ���������� ����       ���������� ���� true     ����������@ ����       ����������@ ����       ���������� ����       ���������� ����       ���������� ����       ���������� ����dec     ���������� ����       ���������� ����       ���������� ����       ���������� ���� true     ���������� ���� true     ���������� ���� true     ���������� ����  false     ���������� ���� true     ���������� ����  false      ���������� ���� true!     ���������� ����  false"     ��������               
                 �� ����       5      ���������� ����       5     ���������� ����       5     ���������� ����       5     ���������� ����       ���������� ����  	     ���������� ����  
     ���������� ����       ���������� ����       ���������� ����       ���������� ���� true     ����������@ ����       ����������@ ����       ���������� ����       ���������� ����       ���������� ����       ���������� ����dec     ���������� ����       ���������� ����       ���������� ����       ���������� ���� true     ���������� ���� true     ���������� ���� true     ���������� ����  false     ���������� ���� true     ���������� ����  false      ���������� ���� true!     ���������� ����  false"     ��������               
                 ��@ ����        ����������@ ����       ���������� ����       ���������� ����       ���������� ����       ���������� ����       ���������� ����       ���������� ����       ���������� ����decade     ���������� ���� true     ���������� ���� true     ���������� ���� true     ���������� ����  false     ��������               
                 �� ����        ���������� ����       ����������@ ����       ����������  ����       ���������� ����       ���������� ����       ���������� ����       ���������� ����       ���������� ����       ���������� ����       ���������� ����       ��������               
                        �� ����dec     ���������� ����     @�@1k     ���������� ����    ��.A1meg     ���������� ����       20     ���������� ����        0     ���������� ����        0     ���������� ���� true	     ���������� ���� true
     ���������� ����      I@50     ���������� ���� true     ���������� ����  false     ��������               
                          / �� ���� x'     ����������     �-���q=1E-12     ���������� @B -C��6?1E-4     ���������� ���� x     ���������� ���� x     ���������� ���� x     ���������� ���� x     ���������� ���� x     ���������� ���� x     ���������� ���� x	     ���������� ���� x!     ���������� ����    �  500
     ���������� ���� x     ���������� ����    �  500     ���������� ���� x$     ���������� ���� x$     ���������� ���� x%     ���������� ���� x"     ����������  ���� x*     ���������� ���� x     ���������� ���� x     ���������� ���� x     ���������� ���� x&     ���������� ���� x     ���������� ���� x     ���������� ���� x     ���������� ���� x+     ���������� ���� x,     ���������� ���� x-     ���������� ���� xg     ���������� ���� xf     ���������� ���� xd     ���������� ���� xe     ���������� ���� xh     ���������� ���� xj     ���������� ���� xi     ���������� ���� xk     ���������� ����    e��A1Gl     ����������             0�     ���������� ����      @5�     ���������� ����      @2.5�     ���������� ����      �?.5�     ���������� ����      @4.5�     ���������� 
   ��&�.>1n�     ���������� 
   ��&�.>1n�     ���������� 
   ��&�.>1n�     ���������� 
   ��&�.>1n�     ��������                                  Ariald        �ڬtd�  ۬t�� ���t    �ڬtd�  ۬t�� ���t ��  COpAnal                         
                        ����                                   �ڬtd�  ۬t�� ���t    �ڬtd�  ۬t�� ���t ��  CDCsweep       
 ����������               
                      ����                                   �ڬtd�  ۬t�� ���t    �ڬtd�  ۬t�� ���t ��  CACsweep        ��������               
                      ����                                  �ڬtd�  ۬t�� ���t    �ڬtd�  ۬t�� ���t �� 
 CTranSweep        ��������               
                      ����                                   �ڬtd�  ۬t�� ���t    �ڬtd�  ۬t�� ���t ��  CACdisto        �����               
                          ����                                  �ڬtd�  ۬t�� ���t    �ڬtd�  ۬t�� ���t ��        �� ����        ���������� ����       ���������� ����       ���������� ����dec     ���������� ����       ��������               
                         ����                                  �ڬtd�  ۬t�� ���t    �ڬtd�  ۬t�� ���t ��        �� ����        ���������� ����       ���������� ����       ���������� ����dec     ���������� ����       ��������               
         �                ����                                  �ڬtd�  ۬t�� ���t    �ڬtd�  ۬t�� ���t ��        �� ����        ���������� ����       ���������� ����       ���������� ����dec     ���������� ����       ��������               
                          ����                                  �ڬtd�  ۬t�� ���t    �ڬtd�  ۬t�� ���t ��        �� ����        ���������� ����       ���������� ����       ���������� ����dec     ���������� ����       ��������               
                         ����                                  �ڬtd�  ۬t�� ���t    �ڬtd�  ۬t�� ���t ��        �� ����        ���������� ����       ���������� ����       ���������� ����dec     ���������� ����       ��������               
         �            	    ����                                  �ڬtd�  ۬t�� ���t    �ڬtd�  ۬t�� ���t ��  CACnoise        ��������               
                   
    ����                                  �ڬtd�  ۬t�� ���t    �ڬtd�  ۬t�� ���t ԃ         ��  ����        ����������  ����       ����������  ����       ���������� ����dec     ���������� ����       ���������� ����       ���������� ����  	     ���������� ����  
     ��������              
                        ����                                  �ڬtd�  ۬t�� ���t    �ڬtd�  ۬t�� ���t ��  CFourier        ����               
         ��                  ����                                   �ڬtd�  ۬t�� ���t    �ڬtd�  ۬t�� ���t ��  CACpz        	 ���������               
                       ����                                   �ڬtd�  ۬t�� ���t    �ڬtd�  ۬t�� ���t ��  CDCtf         �����               
                       ����                                   �ڬtd�  ۬t�� ���t    �ڬtd�  ۬t�� ���t ��  CDCsens         �����������               
                       ����                                   �ڬtd�  ۬t�� ���t    �ڬtd�  ۬t�� ���t                 ����                                   �ڬtd�  ۬t�� ���t    �ڬtd�  ۬t�� ���t ��  CShow         �              
                       ����                                   �ڬtd�  ۬t�� ���t    �ڬtd�  ۬t�� ���t ��  CShowmod         �              
                       ����                                   �ڬtd�  ۬t�� ���t    �ڬtd�  ۬t�� ���t �� 
 CLinearize        ��  ����        ��������               
                      ����                                   �ڬtd�  ۬t�� ���t    �ڬtd�  ۬t�� ���t ��  CParamTranSweep        �������������               
                      ����                                   �ڬtd�  ۬t�� ���t    �ڬtd�  ۬t�� ���t �             ����                                   �ڬtd�  ۬t�� ���t    �ڬtd�  ۬t�� ���t ��  CParamACSweep        Z[\]^_`abcdef               
                      ����                                  �ڬtd�  ۬t�� ���t    �ڬtd�  ۬t�� ���t ��  CMonteCarlo_op        ����������������������                
                             ����                                   �ڬtd�  ۬t�� ���t    �ڬtd�  ۬t�� ���t ��  CMonteCarlo_dc        	
 !               
                      ����                                   �ڬtd�  ۬t�� ���t    �ڬtd�  ۬t�� ���t ��  CMonteCarlo_ac        "#$%&'()*+,-./0123456789:;<=               
                      ����                                  �ڬtd�  ۬t�� ���t    �ڬtd�  ۬t�� ���t ��  CMonteCarlo_tran        >?@ABCDEFGHIJKLMNOPQRSTUVWXY               
                      ����                                   �ڬtd�  ۬t�� ���t    �ڬtd�  ۬t�� ���t ��  CACsens        ghijklmnopq               
                             ����                                  �ڬtd�  ۬t�� ���t    �ڬtd�  ۬t�� ���t ��  CNetworkAnalysis        rstuvwxyz{|               
                      ����                                  �ڬtd�  ۬t�� ���t    �ڬtd�  ۬t�� ���t                 ����                                 >           ��   CDigSimResTemplate                     ��   TDigitalSignal            U1    ���� ����                         �            Q2    ���� ����                         �            Q1    ���� ����                         �            Q0    ���� ����                         �            In1    ���� ����                         �            In2    ���� ����                         �            In3    ���� ����                         �            In4    ���� ����                                  ���       ����  ����:�0�yU>+20.00n���   ����                       Arial����                       Arial����                       Arial                                          ����  ����        0��          ����  ����        0��                     �               ����  �����      1000������          0.000000e+000��    ��������      0.000000e+000��    ��������      0.000000e+000��    ��������   ����                       Arial����                       Arial����                       Arial����                       Arial                        �     �   �  �                     ����  ��    ��������   @  DO14�14 pin small outline package                                                                                                                                                                                                                              ����   ��   CPackageAliasSuperPCBStandardSO14      	�EagleBURR.LBRSO14      	�Orcad SOG.050/14/WG.244/L.350      	�Pads SO14NB      	�	UltiboardL7IC.l55$SO14      	�Eagleburr-brown.lbrSO14             B              @  DO14�14 pin small outline package                                                                                                                                                                                                                              ����   
        A              @  DO14�14 pin small outline package                                                                                                                                                                                                                              ����   	�SuperPCBStandardSO14      	�EagleBURR.LBRSO14      	�Orcad SOG.050/14/WG.244/L.350      	�Pads SO14NB      	�	UltiboardL7IC.l55$SO14      	�Eagleburr-brown.lbrSO14             A              �   DIP-14�14 pin dual in line package                                                                                                                                                                                                                               �     	�SuperPCBStandardDIP14      	�EagleBURR.LBRDIP-14      	�Orcad DIP.100/14/W.300/L.700      	�Pads DIP14      	�	UltiboardUltilib.l55DIP14      	�Eagleburr-brown.lbrDIL14      	�Eagledil.lbrDIL14     	�Eagleanalog-devicesDIL14      	�Eagle74xx-usDIL14      	�Eagle	74ttl-dinDIL14      	�EaglemaximDIL14      	�EagleexarDIL14      	�Eagle
ic-packageDIL14      	�Eagleresistor-dilDIL14      	�EagletexasDIL14      	�Eagle
74ac-logicDIL14              A                                                                                                  �   DIP-14�14 pin dual in line package                                                                                                                                                                                                                               �      !"#$%        B                              �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                   �#     �����  a	    ��     J   J   �      a	J                  2         �                 � � �           u m     ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                   �#     �����  a	    ��     J   J   �      a	J                  2         �                 � � �           u m     ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                   �#     �����  a	    ��     J   J   �      a	J                  2         �                 � � �           u m     ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                   �#     �����  a	    ��     J   J   �      a	J                  2         �                 � � �           u m     ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                   �#     �����  a	    ��     J   J   �      a	J                  2         �                 � � �           u m     ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                   �#     �����  a	    ��     J   J   �      a	J                  2         �                 � � �           u m     ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                   �#     �����  a	    ��     J   J   �      a	J                  2         �                 � � �           u m     ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                   �#     �����  a	    ��     J   J   �      a	J                  2         �                 � � �           u m     ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                   �#     �����  a	    ��     J   J   �      a	J                  2         �                 � � �           u m     ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                   �#     �����  a	    ��     J   J   �      a	J                  2         �                 � � �           u m     ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                   �#     �����  a	    ��     J   J   �      a	J                  2         �                 � � �           u m     ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                   �#     �����  a	    ��     J   J   �      a	J                  2         �                 � � �           u m     ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                   �#     �����  a	    ��     J   J   �      a	J                  2         �                 � � �           u m     ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                   �#     �����  a	    ��     J   J   �      a	J                  2         �                 � � �           u m     ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                   �#     �����  a	    ��     J   J   �      a	J                  2         �                 � � �           u m     ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                   �#     �����  a	    ��     J   J   �      a	J                  2         �                 � � �           u m     ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                   �#     �����  a	    ��     J   J   �      a	J                  2         �                 � � �           u m     ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                   �#     �����  a	    ��     J   J   �      a	J                  2         �                 � � �           u m     ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                   �#     �����  a	    ��     J   J   �      a	J                  2         �                 � � �           u m     ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                   �#     �����  a	    ��     J   J   �      a	J                  2         �                 � � �           u m     ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                   �#     �����  a	    ��     J   J   �      a	J                  2         �                 � � �           u m     ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                   �#     �����  a	    ��     J   J   �      a	J                  2         �                 � � �           u m     ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                   �#     �����  a	    ��     J   J   �      a	J                  2         �                 � � �           u m     ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                   �#     �����  a	    ��     J   J   �      a	J                  2         �                 � � �           u m     ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                   �#     �����  a	    ��     J   J   �      a	J                  2         �                 � � �           u m     ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                   �#     �����  a	    ��     J   J   �      a	J                  2         �                 � � �           u m     ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                   �#     �����  a	    ��     J   J   �      a	J                  2         �                 � � �           u m     ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                   �#     �����  a	    ��     J   J   �      a	J                  2         �                 � � �           u m     ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                   �#     �����  a	    ��     J   J   �      a	J                  2         �                 � � �           u m     ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                   �#     �����  a	    ��     J   J   �      a	J                  2         �                 � � �           u m     ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                               �� 	 CTitleBox                                                      �	                  ?�         �  @                  ���                                                  �  @  A�     <   �  <     ��                                                        A�     |   �  |     ��                                                        A�     �   �  �     ��    � <                                                 A�     �   �  �     ��                                                        E� h      t  4     ��                                                      h      t  4   h      t  4   [title]                                       E� �   H   �  x     ��                                                      �   H   �  x   �   H   �  x   [description]                                       E� P   �   X  �     ��                                                      P   �   X  �   P   �   X  �   [id]                                       E� �   �   �  �     ��                                                      �   �   �  �   �   �   �  �   
[designer]                                       E�      ]   1    ��        	                                                   ]   1       ]   1  Date :       �  4  �  �                  E� p     x  4   	 ��        
                                              p     x  4  p     x  4  [date]                                       E�       U   1    
 ��                                                            U   1         U   1   Title :       �  4  �  �                  E�    L   �   q     ��                                                         L   �   q      L   �   q   Description :       �  �  �   �                  E�    �   8   �     ��                                                         �   8   �      �   8   �   ID :       �  �  8  J                  E�    �   �   �     ��                                                         �   �   �      �   �   �   
Designer :       �  t  p   
                   ()*+,-./023456          1     	title box     Miscellaneous      �?    9 
 ��  CParamSubBehavior    
 ��  ����        ����������  ����       ����������  ����       ����������  ����       ����������  ����       ����������  ����       ����������  ����       ����������  ����       ����������  ����       ����������  ����  	     ��������        9                                      ������   CParamSubModelType�� ����  
   ��  	 CParmDefn            title                E�            description                E�            id                E�            designer                E�            Date :                E�            date                E�            Title :                E�            Description :                E�            ID :                E�            
Designer :                            ����             `         �?�� 	 CGraphDoc�  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                                                                                            2         �                 � � �                   ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                         U1Q2Q1Q0In1In2In3In4                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          1m  0                            100   100                                                           1m  0                            100   100                              1m  0                            100   100                              1m  0                            100   100                                                 
               1m  0                            100   100                            ��   CPartPackage     ��   CPackage@  DO14�14 pin small outline package                                                                                                                                                                                                                              ����   
   R��� T�@  DO14�14 pin small outline package                                                                                                                                                                                                                              ����      R�    T��   DIP-14�14 pin dual in line package                                                                                                                                                                                                                               �      !"#$%   S ��   CMiniPartPin    ����JJ     INJ�      Z�   ����CkCk     INCk�     Z�   ����KK     INK�     Z�   ����RR     INR�     Z�   ����QQ     OUTQ�     Z�   ����Q'Q'     OUTQ'�          ��   CPackagePin 10 RIN 
 BB.Ra� 1 JIN  AJa� 4 KIN  AKa� 8 JIN  BB.Ja� 11 KIN  BB.Ka� 3 QOUT  AA.Qa� 2 Q'OUT  AA.Q'a� 13 RIN  AA.Ra� 5 QOUT  BB.Qa� 6 Q'OUT  BB.Q'a� 9 CkIN 	 BB.Clka� 12 CkIN  AA.ClkJK Flip-Flop w/clear
Flip FlopsGenericC      74107 A74107DA1               DIP1474107D74107D��  CXSpiceBehavior       jkclkresetoutnout ��   CBehPin     j����    �  j����                         ��p�    k����   �  k����                         ��p�    clk����   �  clk����                         ��p�     set����   �  set����                         ��p�    reset����   �  reset����                         ��p�    out����   �  out����                        ��p�    nout����   �  nout����                        ��74107 (XSpice)74107 (XSpice)  8               qrstuvwDigital<   Generic               ����    * time value noutQ'jJkKresetRoutQclkCk CkclkJjKkQ'noutQoutRreset                                                     S Z�    ����JJ     INJ�      Z�   ����CkCk     INCk�     Z�   ����KK     INK�     Z�   ����RR     INR�     Z�   ����QQ     OUTQ�     Z�   ����Q'Q'     OUTQ'�          bcdefghijklmJK Flip-Flop w/clear
Flip FlopsGenericC      74107 A74107DA1               DIP1474107D74107Dn�       jkclkresetoutnout p�     j����    �  j����                         ��p�    k����   �  k����                         ��p�    clk����   �  clk����                         ��p�     set����   �  set����                         ��p�    reset����   �  reset����                         ��p�    out����   �  out����                        ��p�    nout����   �  nout����                        ��74107 (XSpice)74107 (XSpice)  8               ������Digital<   Generic               ����    * time value noutQ'jJkKresetRoutQclkCk CkclkJjKkQ'noutQoutRreset                                                     V Z�    ����JJ     INJ�      Z�   ����CkCk     INCk�     Z�   ����KK     INK�     Z�   ����RR     INR�     Z�   ����QQ     OUTQ�     Z�   ����Q'Q'     OUTQ'�         a� 10 RPassive 
 BB.Ra� 1 JIN  AJa� 4 KIN  AKa� 8 JPAS  BB.Ja� 11 KPAS  BB.Ka� 3 QOUT  AA.Qa� 2 Q'OUT  AA.Q'a� 13 RIN  AA.Ra� 5 QPassive  BB.Qa� 6 Q'PAS  BB.Q'a� 9 CkPassive 	 BB.Clka� 12 CkIN  AA.ClkJK Flip-Flop w/clear
Flip FlopsGenericC      74107 A74107DA2                DIP1474107D74107Dn�       jkclkresetoutnout p�     j����    �  j����                         ��p�    k����   �  k����                         ��p�    clk����   �  clk����                         ��p�     set����   �  set����                         ��p�    reset����   �  reset����                         ��p�    out����   �  out����                        ��p�    nout����   �  nout����                        ��74107 (XSpice)74107 (XSpice)  8               �������Digital<   Generic               ����    * time value noutQ'jJkKresetRoutQclkCk CkclkJjKkQ'noutQoutRreset                                                     X Z�    ����aA     IN1AA  �?  Z�   ����bB     IN1BB  �?  Z�   ����yY     OUT1Y@  �?    #   a� 1 a   A1Aa� 2 b   A1Ba� 3 y   A1Ya� 4 a   B2Aa� 5 b   B2Ba� 6 y   B2Ya� 7  GND  COMGNDa� 8 y   C3Ya� 9 a  	 C3Aa� 10 b  
 C3Ba� 11 y   D4Ya� 12 a   D4Aa� 13 b   D4Ba� 14  VCC  COMVCCXSpice 2input AND gateGatesGeneric=      7408 A74LS08NA3                       DIP1474LS08N74LS08Nn�       aby p� �?  a����    �  a����                        ��p� �?  b����   �  b����                        ��p� �?  y����   �  y����                        ��7408 LS 2-input And7408 LS 2-input And  8               ���Digital<   Generic                       * time value yYaAbB YyAaBb                                Z�    ����AA     INA�      ClockClock                  Z�    ����portport       ��������Output_PortOutput_Port                  Z�    ����portport       ��������Output_PortOutput_Port                  Z�    ����portport       ��������Output_PortOutput_Port                  Z�    ����AA     INA      InputInput                  Z�    ����AA     INA      InputInput                  Z�    ����aA     INaE      Z�   ����bB     INbD     Z�   ����cC     INcF     Z�   ����yY     OUTyC     74ALS11A74ALS11A                                       X Z�    ����aA     IN1AA  �?  Z�   ����bB     IN1BB  �?  Z�   ����yY     OUT1Y@  �?    #   ��������������XSpice 2input AND gateGatesGeneric=      7408 A74LS08NA3                       DIP1474LS08N74LS08Nn�       aby p� �?  a����    �  a����                        ��p� �?  b����   �  b����                        ��p� �?  y����   �  y����                        ��7408 LS 2-input And7408 LS 2-input And  8               ���Digital<   Generic                       * time value yYaAbB YyAaBb                                Z�    ����AA     INA      InputInput                  Z�    ����AA     INA      InputInput                                                         