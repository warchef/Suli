    � B2SPICE zzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzz  
  ��  CPart          @           @                 74107D��  CIntPin    ��  CWire      �       �         @           @                 74107D�    �    	 �    
    �         �  �        �  �              7404D �   �    �       9   ��  	 TModelPin    K����   ����K����                          ��      x��    ��������      x��    ��������      x��    ��������      x��    ��������      x��    ��������      x��    �������� d   :�0�yE>10e-9��    �������� d   :�0�yE>10e-9��    ��������                             ����  ����:�0�yE>10e-9��d         ����  ����:�0�yE>10e-9��d   �      ��   TJKFF_general       JCkKRQQ' �     J����    ����J����                          ��      x��    ��������      x��    ��������      x��    ��������      x��    ��������      x��    ��������      x��    �������� d   :�0�yE>10e-9��    �������� d   :�0�yE>10e-9��    ��������                             ����  ����:�0�yE>10e-9��d         ����  ����:�0�yE>10e-9��d   �     
    �����     ��   d   :�0�yE>10e-9��    �������� d   :�0�yE>10e-9��    ���������    Ck����   ����Ck����                          ��      x��    ��������      x��    ��������      x��    ��������      x��    ��������      x��    ��������      x��    �������� d   :�0�yE>10e-9��    �������� d   :�0�yE>10e-9��    ��������                            ����  ����:�0�yE>10e-9��d         ����  ����:�0�yE>10e-9��d   �     �    �       11 �        ��   TClock       �   �  �      �   �  �              Clock ��  CExtPin    ��  CVertex9   �  @   ��  CSegment   �   `  @              �    �   �  @   �   # �%   �  �   �/   % �    �  �   & �   �#   �      �   ) �          * �   + �   �      ,                    (     '     �0   ' �<    
  �   . �1   �:    
      0 �-   1 �   �
      2 �$   3 �;   �      4                         /     �   / �?   �  �   �4   �=   �      8 �2   9 �
   @      : �)   ; �I   �      <                        7     6                         $         "                    �     A�                 U1     ��   CPin                   ��                                                       �   `   A�� 
 TRectangle     @   �   �                  ����                                             @   �   �   ��  TLine �   `   �   `     ��    �X                                                B� `   @   `   �     ��    8�W                                                B� p   h   x   h     ��    ��W                                                B� x   T   x   h     ��    X                                                B� x   T   �   T     ��    ��W                                                B� �   T   �   h     ��    �W                                                B� �   h   �   h     ��     X                                                B� �   P   �   p      ��    8�W	                                                ��  
 TTextField    P   Z   u    
 ��        
                                                  P   Z   u      P   Z   u   [period]       P    0  �     P   P   t   K� �   `   �   �    	 ��                                                      �   `   �   �   �   `   �   �   ns          @  p  �  �   `   �   x   K�     �����        ��                                                           �����          �����      	[devname]        ����������������    �����      K�        *   @     ��                                                              *   @          *   @   	[refname]          h  �           �   <    J   I   H   G   F M   L N O E   D   C   ?     A      Clock     Miscellaneous      �?      ��   TClockModel     ��  CValue �  I�����z>100n      ��������R� �  I�����j>50n     �������� A �     A����    ����A����                          ��      x��    ��������      x��    ��������      x��    ��������      x��    ��������      x��    ��������      x��    �������� d   :�0�yE>10e-9��    �������� d   :�0�yE>10e-9��    ��������                             ����  ����:�0�yE>10e-9��d         ����  ����:�0�yE>10e-9��d   �      Q   �����         d   :�0�yE>10e-9��    �������� d   :�0�yE>10e-9��    ��������ClockClock              U Digital InstrumentsO   Generic   U1U1           ����  ��    �������� ����  ��    �������� ����  ��    �������� ����  ��    �������� ����  ��    �������� ����  ��    �������� ����  ��    ��������  al      ����Generic             U ��   CPartPin    ����AA      INAA�  ����Digital InstrumentsDigital Clock inputGeneric                                                                              �'                                   11 �       11 �      �         @           @                 74107D�    �    �   \    5 [ �    \    ��   TOutPort       _   @         _   @                 Output_Port^ �    �   �   
   �'   �3   �   
   c �*   d �5   �  �   e �	   �   �  �   �8   �/   `  �   i     h     g         f     �   f �   @  �   �3   l �N   �  �   m         k                         b     �(   b �4   �   
   o                        �   port     �  `	          Q1     >�                   ��                                                           @   port@�         �   `                   ����                                                 �   `   B�     @       @      ��                                                        ��  TEllipse    8       H                  ����
[negative]               ���                       8       H      8       H   K� (   ,   :   Q     ��                                                      (   ,   `   Q   (   ,   `   Q   [value]       X  �	     z
  (   ,   �   T   K�     $       <     ��                                                           $       <       $       <   [port.nbits]      <       ����            �      "Arial                    $       <   K�     ����M         ��                                                           ����M           ����M       	[refname]       @  H	  �  �	      �����       s   q u v w x r      Output_Port     Miscellaneous      �?      ��   TOutPortModel       port � ����port����        port����                                         0��    ��������             0��    ��������             0��    ��������             0��    ��������             0��    ��������             0��    �������� d   :�0�yE>10e-9��    �������� d   :�0�yE>10e-9��    ��������                             ����  ����:�0�yE>10e-9��d         ����  ����:�0�yE>10e-9��d   �     \ z   �����     ��   d   :�0�yE>10e-9��    �������� d   :�0�yE>10e-9��    ��������Output_PortOutput_Port   �            { Digital<   Generic   Q1Q1           ����  ��    �������� ����  ��    �������� ����  ��    �������� ����  ��    �������� ����  ��    �������� ����  ��    �������� ����  ��    ��������          ����       ����  Out V�    ����portport       A X]      Digital Instruments Generic                                                                                                             5  { �    Q����   ����Q����                         �� �  :�0�ye>40ns��    ��������      x��    �������� �   I�����Z>25ns��    �������� �   I�����Z>25ns��    ��������      x��    �������� �   ��&�.Q>16ns��    �������� d   :�0�yE>10e-9��    �������� d   :�0�yE>10e-9��    ��������                            ����  ����:�0�yE>10e-9��d         ����  ����:�0�yE>10e-9��d   �     \ �       JCkKRQQ' �     J����    ����J����                          ��      x��    ��������      x��    ��������      x��    ��������      x��    ��������      x��    ��������      x��    �������� d   :�0�yE>10e-9��    �������� d   :�0�yE>10e-9��    ��������                             ����  ����:�0�yE>10e-9��d         ����  ����:�0�yE>10e-9��d   �      ~   �����     ��   d   :�0�yE>10e-9��    �������� d   :�0�yE>10e-9��    ���������    Ck����   ����Ck����                          ��      x��    ��������      x��    ��������      x��    ��������      x��    ��������      x��    ��������      x��    �������� d   :�0�yE>10e-9��    �������� d   :�0�yE>10e-9��    ��������                            ����  ����:�0�yE>10e-9��d         ����  ����:�0�yE>10e-9��d   �      ~   �����     ��   d   :�0�yE>10e-9��    �������� d   :�0�yE>10e-9��    ���������    K����   ����K����                          ��      x��    ��������      x��    ��������      x��    ��������      x��    ��������      x��    ��������      x��    �������� d   :�0�yE>10e-9��    �������� d   :�0�yE>10e-9��    ��������                             ����  ����:�0�yE>10e-9��d         ����  ����:�0�yE>10e-9��d   �     �    �   �    3 �   �    3 �    �   �
       �   �  p      �   �  p              74ALS11A� �   �    �   �    6 �   �   Z 6 �  �    Q'����   ����Q'����                         �� �  :�0�ye>40ns��    ��������      x��    �������� �   I�����Z>25ns��    �������� �   I�����Z>25ns��    ��������      x��    �������� �   ��&�.Q>16ns��    �������� d   :�0�yE>10e-9��    �������� d   :�0�yE>10e-9��    ��������                           ����  ����:�0�yE>10e-9��d         ����  ����:�0�yE>10e-9��d   �     � ~   �����        d   :�0�yE>10e-9��    �������� d   :�0�yE>10e-9��    ���������    K����   ����K����                          ��      x��    ��������      x��    ��������      x��    ��������      x��    ��������      x��    ��������      x��    �������� d   :�0�yE>10e-9��    �������� d   :�0�yE>10e-9��    ��������                             ����  ����:�0�yE>10e-9��d         ����  ����:�0�yE>10e-9��d   �     � �       JCkKRQQ' �     J����    ����J����                          ��      x��    ��������      x��    ��������      x��    ��������      x��    ��������      x��    ��������      x��    �������� d   :�0�yE>10e-9��    �������� d   :�0�yE>10e-9��    ��������                             ����  ����:�0�yE>10e-9��d         ����  ����:�0�yE>10e-9��d   �     \ �   �����     ��   d   :�0�yE>10e-9��    �������� d   :�0�yE>10e-9��    ���������    Ck����   ����Ck����                          ��      x��    ��������      x��    ��������      x��    ��������      x��    ��������      x��    ��������      x��    �������� d   :�0�yE>10e-9��    �������� d   :�0�yE>10e-9��    ��������                            ����  ����:�0�yE>10e-9��d         ����  ����:�0�yE>10e-9��d   �      �   �����     ��   d   :�0�yE>10e-9��    �������� d   :�0�yE>10e-9��    ��������� �    R����   ����R����                          ��      x��    ��������      x��    ��������      x��    ��������      x��    ��������      x��    ��������      x��    �������� d   :�0�yE>10e-9��    �������� d   :�0�yE>10e-9��    ��������                            ����  ����:�0�yE>10e-9��d         ����  ����:�0�yE>10e-9��d   �     �    �   �    12 �   �   Z 12 �   �    12 �    �    ��   TInPort	       _   @         _   @                 Input� �    �U   �
      �J   �G   `	      �     �     �>   � �B   @      �   �A   @  �   �   �"   @  �   �5   �   @      �6   �@   @  `   �     �     �        �     �     �     �     �     � �=   � �H          �<   �C   �      �7   �D   �      � �"   �   `      �#   �E          �     �     �        �         �     �     �     �   �!   �      �   � �0      `   �         �         �     �                    	        @  �   A   @  @          In1     >�                    ��                                                       �   @   At� �   8   �   H                  ����
[negative]               ���                    �   8   �   H   �   8   �   H   @� t       �   @                   ����A                                      t       �   @   @� t   @   �   `                   ����A                                      t   @   �   `   B� �   @   �   @     ��                                                        @�         �   `                   ����                                                 �   `   B� t       t   `     
 ��                                                      ��  TPolygon                    ��                                                       ��  TPoint�   \       ���   P       ���   P       ���   D       ���   D    `  ���   P       ���   P    `yW    ��                    ��                                                       ���   $       ���   0    `  ���   0        ���   <       ���   <    �  ���   0    �  ���   0    `xW    K� �       �   8    	 ��        	                                               �       �   8   �       �   8   	[A.nbits]      <       ����            �      "Arial                �       �   8   K�    (      M     ��        
                                                 (      M      (      M   [value]       L  �  �  N     (   l   P   K� ��������+   #     ��                                                       ��������+   #   ��������+   #   	[refname]       :  1  �  �  ���������       � �   �   � �   � � � � �   � �      input_general     Miscellaneous      �?      ��   TInPortModel       A �     A����    ����A����                         ��             0��    ��������             0��    ��������             0��    ��������             0��    ��������             0��    ��������             0��    �������� d   :�0�yE>10e-9��    �������� d   :�0�yE>10e-9��    ��������                            ����  ����:�0�yE>10e-9��d         ����  ����:�0�yE>10e-9��d   �     � �   �����         d   :�0�yE>10e-9��    �������� d   :�0�yE>10e-9��    ��������1 Bit Inport1 Bit Inport   �t            � Digital<   Generic   In1In1           ����  ��    �������� ����  ��    �������� ����  ��    �������� ����  ��    �������� ����  ��    �������� ����  ��    �������� ����  ��    ��������  Lo�    ����             In V�    ����AA      INAAQ  ����Digital Instruments Generic                         `   `              `   �  �              `   �             �  `   `          �      12  �    R����   ����R����                          ��      x��    ��������      x��    ��������      x��    ��������      x��    ��������      x��    ��������      x��    �������� d   :�0�yE>10e-9��    �������� d   :�0�yE>10e-9��    ��������                            ����  ����:�0�yE>10e-9��d         ����  ����:�0�yE>10e-9��d   �     � ~   �����     ��   d   :�0�yE>10e-9��    �������� d   :�0�yE>10e-9��    ���������    R����   ����R����                          ��      x��    ��������      x��    ��������      x��    ��������      x��    ��������      x��    ��������      x��    �������� d   :�0�yE>10e-9��    �������� d   :�0�yE>10e-9��    ��������                            ����  ����:�0�yE>10e-9��d         ����  ����:�0�yE>10e-9��d   �     �    �����     ��   d   :�0�yE>10e-9��    �������� d   :�0�yE>10e-9��    ��������� �  12�   �����     ��   d   :�0�yE>10e-9��    �������� d   :�0�yE>10e-9��    ���������    Q����   ����Q����                         �� �  :�0�ye>40ns��    ��������      x��    �������� �   I�����Z>25ns��    �������� �   I�����Z>25ns��    ��������      x��    �������� �   ��&�.Q>16ns��    �������� d   :�0�yE>10e-9��    �������� d   :�0�yE>10e-9��    ��������                            ����  ����:�0�yE>10e-9��d         ����  ����:�0�yE>10e-9��d   �     �    �   �   Z 13 �    �    _�       _   @         _   @                 Output_Port� �    �   @   
   �%   �2   @  �	   �     �     �&   � �   @  �   � �   �   �  �   �   �>   �  �   �     �     �        �                            �   port     @  `	          Q0     >�                   ��                                                           @   port@�         �   `                   ����                                                 �   `   B�     @       @      ��                                                        t�    8       H                  ����
[negative]               ���                       8       H      8       H   K� (   ,   :   Q     ��                                                      (   ,   `   Q   (   ,   `   Q   [value]       �  �	  `  z
  (   ,   �   T   K�     $       <     ��                                                           $       <       $       <   [port.nbits]      <       ����            �      "Arial                    $       <   K�     ����M         ��                                                           ����M           ����M       	[refname]       �  H	  (  �	      �����       �   � � � � � �      Output_Port     Miscellaneous      �?      y�       port � ����port����        port����                                         0��    ��������             0��    ��������             0��    ��������             0��    ��������             0��    ��������             0��    �������� d   :�0�yE>10e-9��    �������� d   :�0�yE>10e-9��    ��������                             ����  ����:�0�yE>10e-9��d         ����  ����:�0�yE>10e-9��d   �     � �   �����     ��   d   :�0�yE>10e-9��    �������� d   :�0�yE>10e-9��    ��������Output_PortOutput_Port   �            � Digital<   Generic   Q0Q0           ����  ��    �������� ����  ��    �������� ����  ��    �������� ����  ��    �������� ����  ��    �������� ����  ��    �������� ����  ��    ��������          ����       ����  Out V�    ����portport       A �>      Digital Instruments Generic                                                                                                             13  � �  13�   �����         d   :�0�yE>10e-9��    �������� d   :�0�yE>10e-9��    ���������    Q'����   ����Q'����                         �� �  :�0�ye>40ns��    ��������      x��    �������� �   I�����Z>25ns��    �������� �   I�����Z>25ns��    ��������      x��    �������� �   ��&�.Q>16ns��    �������� d   :�0�yE>10e-9��    �������� d   :�0�yE>10e-9��    ��������                           ����  ����:�0�yE>10e-9��d         ����  ����:�0�yE>10e-9��d   �     �	    �   �  	 Z 14 �   �  	 � 14  � �    C����   ����C����                          ��      x��    ��������      x��    ��������      x��    ��������      x��    ��������      x��    ��������      x��    �������� d   :�0�yE>10e-9��    �������� d   :�0�yE>10e-9��    ��������                             ����  ����:�0�yE>10e-9��d         ����  ����:�0�yE>10e-9��d   �     � ��   TAnd       ABCY �     A����    ����A����                          ��      x��    ��������      x��    ��������      x��    ��������      x��    ��������      x��    ��������      x��    �������� d   :�0�yE>10e-9��    �������� d   :�0�yE>10e-9��    ��������                             ����  ����:�0�yE>10e-9��d         ����  ����:�0�yE>10e-9��d   �     � �   �����     ��   d   :�0�yE>10e-9��    �������� d   :�0�yE>10e-9��    ���������    B����   ����B����                          ��      x��    ��������      x��    ��������      x��    ��������      x��    ��������      x��    ��������      x��    �������� d   :�0�yE>10e-9��    �������� d   :�0�yE>10e-9��    ��������                             ����  ����:�0�yE>10e-9��d         ����  ����:�0�yE>10e-9��d   �     � �   �����     ��   d   :�0�yE>10e-9��    �������� d   :�0�yE>10e-9��    ��������� �    Y����   ����Y����                         �� d   :�0�yE>10ns��    ��������    ��&�.!>2ns��    ��������      x��    �������� �   �?Y��K>13ns��    ��������    ��&�.!>2ns��    ��������      x��    �������� d   :�0�yE>10e-9��    �������� d   :�0�yE>10e-9��    ��������                            ����  ����:�0�yE>10e-9��d         ����  ����:�0�yE>10e-9��d   �     
 �   �����        d   :�0�yE>10e-9��    �������� d   :�0�yE>10e-9��    ��������11A/3 ALS 3-input And11A/3 ALS 3-input And  D �t            � � � � Digital<   Motorola   U3U3           ���� x��    �������� ���� x��    �������� @ �h㈵��>20u��    �������� ����-C��6�-.1m��    �������� ���-C��6:�-.4m��    ��������  ������Mb�?8m��    �������� @]� ��_�LU?1.3m��    ��������         ����ALS      �����     ��   d   :�0�yE>10e-9��    �������� d   :�0�yE>10e-9��    ��������	 14�   �����        d   :�0�yE>10e-9��    �������� d   :�0�yE>10e-9��    ��������107 JK FF w/clear107 JK FF w/clear   �            � � � � � � Digital<   Generic   A3A3           ���� x��    �������� ���� x��    �������� �'	 hUMu?60u��    �������� ʑ�b2U0*�c�-2.4m��    �������� ���-C��6:�-.4m��    ��������  h�	����Mb�?16m��    ��������  ��{�G�z�?10m��    ��������          ����Standard TTL                 0��    �������� ����    �sA20meg��    �������� 6  ��创�`>31n��    ��������             0��    ��������  �����     ��   d   :�0�yE>10e-9��    �������� d   :�0�yE>10e-9��    ���������  6  � 6 � �   
    � 7 �    �'       	   �?   � �J      �
   � �A   �K   �  �
   �@   �*   �  �   �   �   �  `   �   �   �  `   �
   �   �  `                               �   �      �   �   	�    �  �   
                         �     �     �                
           �  yC  �   �M   �   	   �   �(   �   	           �    �-       	   �   �.      `   �   �   @  `              �   �$   �  `                                  
      �  �  bD  �   �L   �  `	   �D   �Q   �  `	           �E   �P   �	  `	   �C   �O   �	  `   �B   �	   �
  `   �   !�1   @  `   "                     �    �   `	  `   �!   �    	  `   &    %    $                              
       �  �  aE  �   �)   �  �   �F   �T   �  �   * 	   )    �I   )�R   �  �   �G   -�S   �  `   �H   �   �  `   0 	      /    . 	       , 	        	  
      �     cF      �         U3     >�                    ��                                                           �   y>�                   ��                                                      �   �   b>�                   ��                                                      �   �   a>�                   ��                                                      �   `   cB� �   �   �   �     ��     ~�                                                ��   TArc ����p   d   �                                                                  P   �   �      P   �   �   \   P      �           B� �   �   \   �    
 ��    h                                                  7� �����   d      	                                                              0   �   �      0   �   �      �   \   �           B� �   P   \   P     ��    ��                                                B�     �       �     ��    {  	                                                B� �   �   �   �     ��    (��
                                                B� �   `   �   `     ��       �                                                B� �   �   �   P     ��    ��                                                K�         *   H     ��                                                               *   H           *   H   	[refname]          �  �  �          �   D   K�     �����         ��                                                           �����           �����       	[devname]        ����������������    �����        25  3?4>  =  <  ;@A  :  9  8  6   AND 3    
AND 3 IEEEMiscellaneous      �?    D  �   U V�    ����aA      INAaz	  ����V�   ����bB      INAb{	  ����V�   ����cC      INAc|	  ����V�   ����yY      OUTAy}	  ����Gatestriple 3-input AND gatesGeneric               3  � �    Q'����   ����Q'����                         �� �  :�0�ye>40ns��    ��������      x��    �������� �   I�����Z>25ns��    �������� �   I�����Z>25ns��    ��������      x��    �������� �   ��&�.Q>16ns��    �������� d   :�0�yE>10e-9��    �������� d   :�0�yE>10e-9��    ��������                           ����  ����:�0�yE>10e-9��d         ����  ����:�0�yE>10e-9��d   �     �    �����        d   :�0�yE>10e-9��    �������� d   :�0�yE>10e-9��    ���������  3~   �����     ��   d   :�0�yE>10e-9��    �������� d   :�0�yE>10e-9��    ��������� } � 107 JK FF w/clear107 JK FF w/clear   �             � � � } � Digital<   Generic   A2A2           ���� x��    �������� ���� x��    �������� �'	 hUMu?60u��    �������� ʑ�b2U0*�c�-2.4m��    �������� ���-C��6:�-.4m��    ��������  h�	����Mb�?16m��    ��������  ��{�G�z�?10m��    ��������          ����Standard TTL                 0��    �������� ����    �sA20meg��    �������� 6  ��创�`>31n��    ��������             0��    ��������  �����         d   :�0�yE>10e-9��    �������� d   :�0�yE>10e-9��    ���������  5   Z 5 Y � � � � �    l        �  J�  �   ;       �  Ck�  �         @  K�  �   �         R�  �   �   @  �  Q�  �   1  @  @  Q'�   @   
          A3     >�                    ��                                                           �   J>�                   ��                                                          �   Ck>�                   ��                                                          �   K>�                   ��                                                      `      R>�                   ��                                                      �   �   Q>�                   ��                                                      �   �   Q'@�     `   �   �                  ����                                             `   �   �   B�     �       �     ��                                                        B�     �       �     ��                                                        B�     �       �    	 ��        	                                                B� `   �   `       
 ��    ����
                                                B� �   �   �   �     ��    ����                                                B� �   �   �   �     ��    ����                                                B� �   x   �   �     ��    ����                                                B� �   x   �   x     ��    ����                                                t� X   �   h   �                  �                                           X   �   h   �   X   �   h   �   B� �   �   �   �     ��    ����                                                B� �   �   �   �     ��    ����                                                t� �   �   �   �                  �                                           �   �   �   �   �   �   �   �   K�     0   b   X     ��                                                           0   b   X       0   b   X   	[refname]       �  �
  h  P      0   �   T   K� (   p   0   �     ��                                                      (   p   0   �   (   p   0   �   j       �  p  �    (   p   p   �   K� (   �   P   �     ��                                                      (   �   P   �   (   �   P   �   clk       �  �  0  f  (   �   p   �   K� (   �   8   �     ��                                                      (   �   8   �   (   �   8   �   k       �  0  �  �  (   �   p   �   K�        �   0     ��                                                              �   0          �   0   	[devname]        ����������������       �   0    MNOPQRSTUVWXYabc      [  ]^dZ_`  \     74107 JK FF w/clear    74107 JK FF w/clear IEEEMiscellaneous      �?      �   A V�    ����JJ      INAJ�>  ����V�   ����CkCk      INACk�>  ����V�   ����KK      INAK�>  ����V�   ����RR      INAR�>  ����V�   ����QQ      OUTAQ    ����V�   ����Q'Q'      OUTAQ'��/A����V�    ����JJ      INBJ    ����V�   ����CkCk      INBCk�>  ����V�   ����KK      INBK��������V�   ����RR      INBR�>  ����V�   ����QQ      OUTBQ�>  ����V�   ����Q'Q'      OUTBQ'�>  ����
Flip FlopsJK Flip-Flop w/clearGenericDO14              11  �  � U  11   �����     ��   d   :�0�yE>10e-9��    �������� d   :�0�yE>10e-9��    �������� � �    Q����   ����Q����                         �� �  :�0�ye>40ns��    ��������      x��    �������� �   I�����Z>25ns��    �������� �   I�����Z>25ns��    ��������      x��    �������� �   ��&�.Q>16ns��    �������� d   :�0�yE>10e-9��    �������� d   :�0�yE>10e-9��    ��������                            ����  ����:�0�yE>10e-9��d         ����  ����:�0�yE>10e-9��d   �         �����         d   :�0�yE>10e-9��    �������� d   :�0�yE>10e-9��    ��������F107 JK FF w/clear107 JK FF w/clear   �t               � qFDigital<   Generic   A1A1           ���� x��    �������� ���� x��    �������� �'	 hUMu?60u��    �������� ʑ�b2U0*�c�-2.4m��    �������� ���-C��6:�-.4m��    ��������  h�	����Mb�?16m��    ��������  ��{�G�z�?10m��    ��������          ����Standard TTL                 0��    �������� ����    �sA20meg��    �������� 6  ��创�`>31n��    ��������             0��    ��������  �����     ��   d   :�0�yE>10e-9��    �������� d   :�0�yE>10e-9��    ���������    Y����   ����Y����                         �� �   ,i�)+P>15ns��    ��������      x��    �������� d   :�0�yE>10ns��    �������� �   ,i�)+P>15ns��    ��������      x��    �������� Z   h�+e�SC>9ns��    �������� d   :�0�yE>10e-9��    �������� d   :�0�yE>10e-9��    ��������                           ����  ����:�0�yE>10e-9��d         ����  ����:�0�yE>10e-9��d   �      �       InY �     In����    ����In����                          ��      x��    ��������      x��    ��������      x��    ��������      x��    ��������      x��    ��������      x��    �������� d   :�0�yE>10e-9��    �������� d   :�0�yE>10e-9��    ��������                             ����  ����:�0�yE>10e-9��d         ����  ����:�0�yE>10e-9��d   �     
 s  �����     ��   d   :�0�yE>10e-9��    �������� d   :�0�yE>10e-9��    ��������r04/6 LS Inverter04/6 LS Inverter =               trDigital<   Generic   A4A4           ���� x��    �������� ���� x��    �������� @ �h㈵��>20u��    �������� ���-C��6:�-.4m��    �������� ���-C��6:�-.4m��    ��������  ������Mb�?8m��    ��������  6nb2U0*�c?2.4m��    ��������  4�    ����LS      �����         d   :�0�yE>10e-9��    �������� d   :�0�yE>10e-9��    �������� 9   9 �           �  in�  �   �   `  `   �   �,      `   x    w    �   w�      `   z�   {�&   �  `   |                            �  �  out�   �  �
          A4     >�                   ��                                                           �   in>�                   ��                                                      �   �   outt� l   t   �   �                   ���                                          l   t   �   �   l   t   �   �   B� �   �   �   �     ��                                                        B�     �   ,   �     ��                                                        �� ����    ����      ��                                                         ��,   \    �"���,   �    G   ��l   �    �%y@��,   \    S       K� ����   �   0     ��                                                       ����   �   0   ����   �   0   	[devname]        ��������������������   �   0   K� ����0   >   X     ��                                                       ����0   >   X   ����0   >   X   	[refname]       t  p  <    ����0   �   T   	 �  ~�����     Inverter    Inverter IEEEMiscellaneous      �?    =  s  A V�    ����inIn      PASA1AW]  ����V�   ����outY      PASA1YV]  ����V�    ����inIn      PASB1AU]  ����V�   ����outY      PASB1YT]  ����V�    ����inIn      PASC1AS]  ����V�   ����outY      PASC1YR]  ����V�    ����inIn      PASD1AQ]  ����V�   ����outY      PASD1YP]  ����V�    ����inIn      PASE1AO]  ����V�   ����outY      PASE1Y    ����V�    ����inIn      PASF1A    ����V�   ����outY      PASF1Y    ����Gatesdigital one-bit-wide inverterGenericDO14              7 �   t�  7    7 X  �  � �    	       �  J�  �   +       �  Ck�  �   {      @  K�  �   �         R�  �   �   `	  �   �   �+   �  �   �     �    �;   ��8    
  �   �.   �6    
   
   �+   ��   �
   
   ��,   ��7   @   
   �                      �     �    ��:   ��   �
  �   ��9   ��F   @  �   �                                          @  �  Q�  �   %  @  @  Q'�       
          A1     >�                    ��                                                           �   J>�                   ��                                                          �   Ck>�                   ��                                                          �   K>�                   ��                                                      `      R>�                   ��                                                      �   �   Q>�                   ��                                                      �   �   Q'@�     `   �   �                  ����                                             `   �   �   B�     �       �     ��                                                        B�     �       �     ��                                                        B�     �       �    	 ��        	                                                B� `   �   `       
 ��        
                                                B� �   �   �   �     ��                                                        B� �   �   �   �     ��    ����                                                B� �   x   �   �     ��    ����                                                B� �   x   �   x     ��                                                        t� X   �   h   �                  �                                           X   �   h   �   X   �   h   �   B� �   �   �   �     ��                                                        B� �   �   �   �     ��                                                        t� �   �   �   �                  �                                           �   �   �   �   �   �   �   �   K�     0   b   X     ��                                                           0   b   X       0   b   X   	[refname]       �  �
  H  P      0   �   T   K� (   p   0   �     ��                                                      (   p   0   �   (   p   0   �   j       �  p  �    (   p   p   �   K� (   �   P   �     ��                                                      (   �   P   �   (   �   P   �   clk       �  �    f  (   �   p   �   K� (   �   8   �     ��                                                      (   �   8   �   (   �   8   �   k       �  0  �  �  (   �   p   �   K�        �   0     ��                                                              �   0          �   0   	[devname]        ����������������       �   0    ����������������      �  ������  �0     74107 JK FF w/clear    74107 JK FF w/clear IEEEMiscellaneous      �?         A V�    ����JJ      INAJyE>����V�   ����CkCk      INACkE>1����V�   ����KK      INAK    ����V�   ����RR      INAR�<�����V�   ����QQ      OUTAQ   �����V�   ����Q'Q'      OUTAQ'�>  ����V�    ����JJ      INBJ�>  ����V�   ����CkCk      INBCk�>  ����V�   ����KK      INBK�>  ����V�   ����RR      INBR��������V�   ����QQ      OUTBQ�>  ����V�   ����Q'Q'      OUTBQ'�>  ����
Flip FlopsJK Flip-Flop w/clearGenericDO14              1 �         _�       _   @         _   @                 Output_Port��    �       �   port     �
  `	          Q2     >�                   ��                                                           @   port@�         �   `                   ����                                                 �   `   B�     @       @      ��                                                        t�    8       H                  ����
[negative]               ���                       8       H      8       H   K� (   ,   :   Q     ��                                                      (   ,   `   Q   (   ,   `   Q   [value]       �
  �	  �  z
  (   ,   �   T   K�     $       <     ��                                                           $       <       $       <   [port.nbits]      <       ����            �      "Arial                    $       <   K�     ����M         ��                                                           ����M           ����M       	[refname]       �
  H	  h  �	      �����       �  ������     Output_Port     Miscellaneous      �?      y�       port � ����port����        port����                                         0��    ��������             0��    ��������             0��    ��������             0��    ��������             0��    ��������             0��    �������� d   :�0�yE>10e-9��    �������� d   :�0�yE>10e-9��    ��������                             ����  ����:�0�yE>10e-9��d         ����  ����:�0�yE>10e-9��d   �      �  �����     ��   d   :�0�yE>10e-9��    �������� d   :�0�yE>10e-9��    ��������Output_PortOutput_Port                 �Digital<   Generic   Q2Q2           ����  ��    �������� ����  ��    �������� ����  ��    �������� ����  ��    �������� ����  ��    �������� ����  ��    �������� ����  ��    ��������          ����       ����  Out V�    ����portport       A ����    Digital Instruments Generic                                                                                                             1  � q  1  �� 1  � � ] � �    �       �  J�  �   3       �  Ck�  �   !      @  K�  �   �         R�  �   h   @  �  Q�  �     @  @  Q'�   �
   
          A2     >�                    ��                                                           �   J>�                   ��                                                          �   Ck>�                   ��                                                          �   K>�                   ��                                                      `      R>�                   ��                                                      �   �   Q>�                   ��                                                      �   �   Q'@�     `   �   �                  ����                                             `   �   �   B�     �       �     ��                                                        B�     �       �     ��                                                        B�     �       �    	 ��        	                                                B� `   �   `       
 ��    ���
                                                B� �   �   �   �     ��                                                        B� �   �   �   �     ��                                                        B� �   x   �   �     ��                                                        B� �   x   �   x     ��                                                        t� X   �   h   �                  �                                           X   �   h   �   X   �   h   �   B� �   �   �   �     ��    ���                                                B� �   �   �   �     ��                                                        t� �   �   �   �                  �                                           �   �   �   �   �   �   �   �   K�     0   b   X     ��                                                           0   b   X       0   b   X   	[refname]       �
  �
  �  P      0   �   T   K� (   p   0   �     ��                                                      (   p   0   �   (   p   0   �   j       �
  p      (   p   p   �   K� (   �   P   �     ��                                                      (   �   P   �   (   �   P   �   clk       �
  �  p  f  (   �   p   �   K� (   �   8   �     ��                                                      (   �   8   �   (   �   8   �   k       �
  0  (  �  (   �   p   �   K�        �   0     ��                                                              �   0          �   0   	[devname]        ����������������       �   0    ����������������      �  ������  ��     74107 JK FF w/clear    74107 JK FF w/clear IEEEMiscellaneous      �?      ~   A V�    ����JJ      INAJ    ����V�   ����CkCk      INACk   ����V�   ����KK      INAK 5����V�   ����RR      INAR   ����V�   ����QQ      OUTAQ  x����V�   ����Q'Q'      OUTAQ'0e-9����V�    ����JJ      INBJ10e-����V�   ����CkCk      INBCk J�����V�   ����KK      INBK   ����V�   ����RR      INBR d ����V�   ����QQ      OUTBQ �������V�   ����Q'Q'      OUTBQ'yE>����
Flip FlopsJK Flip-Flop w/clearGenericDO14              Z   �` �   � � 
 
 
   � � \ � 
  � � K J K 
�   �                �   �               k g �   � ( 6 , * " |  � z� $ � x� �"$&� � 4 � � c o < e ��2 �& . 0 : m 8 � � � i ���� � � �  �  *.0,� V U V ' - � �h %� !; 	l ! 3 '1�w{� + �b � � #   � � ) % }� )�yj � #� d p f ��� 1 5 / 9 � 7 � � � � � � �� � = � � n -/+�              
 R�@ ����        ��������R�             0     ��������R� ����      @5     ��������R�  ʚ;�������?.1     ��������R�@ ����       ��������R� ����       ��������R� ����       ��������R� ����       ��������R� ���� true
     ��������R� ����  false     ��������               
                  R� ����        ��������R� ����       ��������R�  ����       ��������R�@ ����       ��������R�@ ����       ��������               
                  R� ����        ��������R� ����       ��������R�@ ����       ��������R�  ����       ��������R� ����       ��������R� ����       ��������R� ����       ��������R� ����       ��������R� ����       ��������R� ����       ��������R� ����       ��������               
                 R� ����dec     ��������R� ����     @�@1k     ��������R� ����    ��.A1meg     ��������R� ����       20     ��������R� ���� true     ��������R� ���� true     ��������R� ���� true	     ��������R� ����  false
     ��������               
                 R�  ����        ��������R�  ����       ��������R�  ����       ��������R� ����dec     ��������R� ����       ��������R� ����       ��������R� ����  	     ��������R� ����  
     ��������               
                  	 R� ����        ��������R� ����       ��������R� ����       ��������R� ����       ��������R� ����       ��������R� ����       ��������R� ����       ��������R� ����       ��������R� ����       ��������               
                 R� ����        ��������R� ����       ��������R� ����       ��������R� ����dec     ��������R� ����       ��������               
                     R�             0      ��������R� ��� ����MbP?1m     ��������R� �� �h㈵��>10u     ��������R� '  ���ư>1u     ��������R� ���� true     ��������R� ����  false     ��������R� ���� true     ��������R� ����  false     ��������               
                 R� ����     @�@1K      ��������R�  ����       ��������R�  ����       ��������R�  ����       ��������               
         ��              R�  ����        ��������              
                  R�  ����        ��������              
                                  
                 R�@ ����        ��������R�@ ����       ��������R� ����       ��������R� ����       ��������R� ����       ��������R� ����       ��������R� ����       ��������R� ����       ��������R� ����       ��������R� ���� true	     ��������R� ����  false
     ��������R� ���� true     ��������R� ����  false     ��������               
                 R� ����       5      ��������R� ����       5     ��������R� ����       5     ��������R� ����       5     ��������R� ����       ��������R� ����  	     ��������R� ����  
     ��������R� ����       ��������R� ����       ��������R� ����       ��������R� ���� true     ��������R�@ ����       ��������R�@ ����       ��������R� ����       ��������R� ����       ��������R� ����       ��������R� ����dec     ��������R� ����       ��������R� ����       ��������R� ����       ��������R� ���� true     ��������R� ���� true     ��������R� ���� true     ��������R� ����  false     ��������R� ���� true     ��������R� ����  false      ��������R� ���� true!     ��������R� ����  false"     ��������               
                        R� ����       5      ��������R� ����       5     ��������R� ����       5     ��������R� ����       5     ��������R� ����       ��������R� ����  	     ��������R� ����  
     ��������R� ����       ��������R� ����       ��������R� ����       ��������R� ���� true     ��������R�@ ����       ��������R�@ ����       ��������R� ����       ��������R� ����       ��������R� ����       ��������R� ����dec     ��������R� ����       ��������R� ����       ��������R� ����       ��������R� ���� true     ��������R� ���� true     ��������R� ���� true     ��������R� ����  false     ��������R� ���� true     ��������R� ����  false      ��������R� ���� true!     ��������R� ����  false"     ��������               
                 R� ����       5      ��������R� ����       5     ��������R� ����       5     ��������R� ����       5     ��������R� ����       ��������R� ����  	     ��������R� ����  
     ��������R� ����       ��������R� ����       ��������R� ����       ��������R� ���� true     ��������R�@ ����       ��������R�@ ����       ��������R� ����       ��������R� ����       ��������R� ����       ��������R� ����dec     ��������R� ����       ��������R� ����       ��������R� ����       ��������R� ���� true     ��������R� ���� true     ��������R� ���� true     ��������R� ����  false     ��������R� ���� true     ��������R� ����  false      ��������R� ���� true!     ��������R� ����  false"     ��������               
                 R� ����       5      ��������R� ����       5     ��������R� ����       5     ��������R� ����       5     ��������R� ����       ��������R� ����  	     ��������R� ����  
     ��������R� ����       ��������R� ����       ��������R� ����       ��������R� ���� true     ��������R�@ ����       ��������R�@ ����       ��������R� ����       ��������R� ����       ��������R� ����       ��������R� ����dec     ��������R� ����       ��������R� ����       ��������R� ����       ��������R� ���� true     ��������R� ���� true     ��������R� ���� true     ��������R� ����  false     ��������R� ���� true     ��������R� ����  false      ��������R� ���� true!     ��������R� ����  false"     ��������               
                 R�@ ����        ��������R�@ ����       ��������R� ����       ��������R� ����       ��������R� ����       ��������R� ����       ��������R� ����       ��������R� ����       ��������R� ����decade     ��������R� ���� true     ��������R� ���� true     ��������R� ���� true     ��������R� ����  false     ��������               
                 R� ����        ��������R� ����       ��������R�@ ����       ��������R�  ����       ��������R� ����       ��������R� ����       ��������R� ����       ��������R� ����       ��������R� ����       ��������R� ����       ��������R� ����       ��������               
                        R� ����dec     ��������R� ����     @�@1k     ��������R� ����    ��.A1meg     ��������R� ����       20     ��������R� ����        0     ��������R� ����        0     ��������R� ���� true	     ��������R� ���� true
     ��������R� ����      I@50     ��������R� ���� true     ��������R� ����  false     ��������               
                          / R� ���� x'     ��������R�     �-���q=1E-12     ��������R� @B -C��6?1E-4     ��������R� ���� x     ��������R� ���� x     ��������R� ���� x     ��������R� ���� x     ��������R� ���� x     ��������R� ���� x     ��������R� ���� x	     ��������R� ���� x!     ��������R� ����    �  500
     ��������R� ���� x     ��������R� ����    �  500     ��������R� ���� x$     ��������R� ���� x$     ��������R� ���� x%     ��������R� ���� x"     ��������R�  ���� x*     ��������R� ���� x     ��������R� ���� x     ��������R� ���� x     ��������R� ���� x&     ��������R� ���� x     ��������R� ���� x     ��������R� ���� x     ��������R� ���� x+     ��������R� ���� x,     ��������R� ���� x-     ��������R� ���� xg     ��������R� ���� xf     ��������R� ���� xd     ��������R� ���� xe     ��������R� ���� xh     ��������R� ���� xj     ��������R� ���� xi     ��������R� ���� xk     ��������R� ����    e��A1Gl     ��������R�             0�     ��������R� ����      @5�     ��������R� ����      @2.5�     ��������R� ����      �?.5�     ��������R� ����      @4.5�     ��������R� 
   ��&�.>1n�     ��������R� 
   ��&�.>1n�     ��������R� 
   ��&�.>1n�     ��������R� 
   ��&�.>1n�     ��������                                  Ariald        �ڬt�$k\�  ۬t� ���t    �ڬt�$k\�  ۬t� ���t ��  COpAnal                         
                        ����                                   �ڬt�$k\�  ۬t� ���t    �ڬt�$k\�  ۬t� ���t ��  CDCsweep       
 	
               
                      ����                                   �ڬt�$k\�  ۬t� ���t    �ڬt�$k\�  ۬t� ���t ��  CACsweep        #$%&'()*               
                      ����                                  �ڬt�$k\�  ۬t� ���t    �ڬt�$k\�  ۬t� ���t �� 
 CTranSweep        ABCDEFGH               
                      ����                                   �ڬt�$k\�  ۬t� ���t    �ڬt�$k\�  ۬t� ���t ��  CACdisto        <=>?@               
                          ����                                  �ڬt�$k\�  ۬t� ���t    �ڬt�$k\�  ۬t� ���t &�        R� ����        ��������R� ����       ��������R� ����       ��������R� ����dec     ��������R� ����       ��������               
         �                ����                                  �ڬt�$k\�  ۬t� ���t    �ڬt�$k\�  ۬t� ���t &�        R� ����        ��������R� ����       ��������R� ����       ��������R� ����dec     ��������R� ����       ��������               
                         ����                                  �ڬt�$k\�  ۬t� ���t    �ڬt�$k\�  ۬t� ���t &�        R� ����        ��������R� ����       ��������R� ����       ��������R� ����dec     ��������R� ����       ��������               
                          ����                                  �ڬt�$k\�  ۬t� ���t    �ڬt�$k\�  ۬t� ���t &�        R� ����        ��������R� ����       ��������R� ����       ��������R� ����dec     ��������R� ����       ��������               
         �                ����                                  �ڬt�$k\�  ۬t� ���t    �ڬt�$k\�  ۬t� ���t &�        R� ����        ��������R� ����       ��������R� ����       ��������R� ����dec     ��������R� ����       ��������               
                     	    ����                                  �ڬt�$k\�  ۬t� ���t    �ڬt�$k\�  ۬t� ���t ��  CACnoise        +,-./012               
                   
    ����                                  �ڬt�$k\�  ۬t� ���t    �ڬt�$k\�  ۬t� ���t F�         R�  ����        ��������R�  ����       ��������R�  ����       ��������R� ����dec     ��������R� ����       ��������R� ����       ��������R� ����  	     ��������R� ����  
     ��������              
                        ����                                  �ڬt�$k\�  ۬t� ���t    �ڬt�$k\�  ۬t� ���t ��  CFourier        IJKL               
         ��                  ����                                   �ڬt�$k\�  ۬t� ���t    �ڬt�$k\�  ۬t� ���t ��  CACpz        	 3456789:;               
                       ����                                   �ڬt�$k\�  ۬t� ���t    �ڬt�$k\�  ۬t� ���t ��  CDCtf                        
                       ����                                   �ڬt�$k\�  ۬t� ���t    �ڬt�$k\�  ۬t� ���t ��  CDCsens          !"               
                       ����                                   �ڬt�$k\�  ۬t� ���t    �ڬt�$k\�  ۬t� ���t                 ����                                   �ڬt�$k\�  ۬t� ���t    �ڬt�$k\�  ۬t� ���t ��  CShow         M              
                       ����                                   �ڬt�$k\�  ۬t� ���t    �ڬt�$k\�  ۬t� ���t ��  CShowmod         N              
                       ����                                   �ڬt�$k\�  ۬t� ���t    �ڬt�$k\�  ۬t� ���t �� 
 CLinearize        R�  ����        ��������               
                      ����                                   �ڬt�$k\�  ۬t� ���t    �ڬt�$k\�  ۬t� ���t ��  CParamTranSweep        OPQRSTUVWXYZ[               
                      ����                                   �ڬt�$k\�  ۬t� ���t    �ڬt�$k\�  ۬t� ���t !             ����                                   �ڬt�$k\�  ۬t� ���t    �ڬt�$k\�  ۬t� ���t ��  CParamACSweep        �������������               
                      ����                                  �ڬt�$k\�  ۬t� ���t    �ڬt�$k\�  ۬t� ���t ��  CMonteCarlo_op        \]^_`abcdefghijklmnopqrstuvw               
                             ����                                   �ڬt�$k\�  ۬t� ���t    �ڬt�$k\�  ۬t� ���t ��  CMonteCarlo_dc        xyz{|}~��������������������               
                      ����                                   �ڬt�$k\�  ۬t� ���t    �ڬt�$k\�  ۬t� ���t ��  CMonteCarlo_ac        ����������������������������               
                      ����                                  �ڬt�$k\�  ۬t� ���t    �ڬt�$k\�  ۬t� ���t ��  CMonteCarlo_tran        ����������������������������               
                      ����                                   �ڬt�$k\�  ۬t� ���t    �ڬt�$k\�  ۬t� ���t ��  CACsens        �����������               
                             ����                                  �ڬt�$k\�  ۬t� ���t    �ڬt�$k\�  ۬t� ���t ��  CNetworkAnalysis        �����������               
                      ����                                  �ڬt�$k\�  ۬t� ���t    �ڬt�$k\�  ۬t� ���t                 ����                                 >           ��   CDigSimResTemplate    
           ��   TDigitalSignal            U1    ���� ����                        r�            Q2    ���� ����                        r�            Q1    ���� ����                        r�            Q0    ���� ����                        r�            In1    ���� ����                                  ���       ����  ����:�0�yU>+20.00n���   ����                       Arial����                       Arial����                       Arial                                          ����  ����        0��          ����  ����        0��                     �               ����  �����      1000������          0.000000e+000��    ��������      0.000000e+000��    ��������      0.000000e+000��    ��������   ����                       Arial����                       Arial����                       Arial����                       Arial                        �     �   �  �                     ����  ��    ��������   @  DO14�14 pin small outline package                                                                                                                                                                                                                              ����   ��   CPackageAliasSuperPCBStandardSO14      x�EagleBURR.LBRSO14      x�Orcad SOG.050/14/WG.244/L.350      x�Pads SO14NB      x�	UltiboardL7IC.l55$SO14      x�Eagleburr-brown.lbrSO14             B              @  DO14�14 pin small outline package                                                                                                                                                                                                                              ����   yz{|}~        A              @  DO14�14 pin small outline package                                                                                                                                                                                                                              ����   x�SuperPCBStandardSO14      x�EagleBURR.LBRSO14      x�Orcad SOG.050/14/WG.244/L.350      x�Pads SO14NB      x�	UltiboardL7IC.l55$SO14      x�Eagleburr-brown.lbrSO14             A              @  DO14�14 pin small outline package                                                                                                                                                                                                                              ����   x�SuperPCBStandardSO14      x�EagleBURR.LBRSO14      x�Orcad SOG.050/14/WG.244/L.350      x�Pads SO14NB      x�	UltiboardL7IC.l55$SO14      x�Eagleburr-brown.lbrSO14             A                                                                                  �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                   ��$     ����X� 06`	     �     N   N   n�     06`	N                  2         �                 � � �           u m     ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                   ��$     ����X� 06`	     �     N   N   n�     06`	N                  2         �                 � � �           u m     ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                   ��$     ����X� 06`	     �     N   N   n�     06`	N                  2         �                 � � �           u m     ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                   ��$     ����X� 06`	     �     N   N   n�     06`	N                  2         �                 � � �           u m     ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                   ��$     ����X� 06`	     �     N   N   n�     06`	N                  2         �                 � � �           u m     ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                   ��$     ����X� 06`	     �     N   N   n�     06`	N                  2         �                 � � �           u m     ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                   ��$     ����X� 06`	     �     N   N   n�     06`	N                  2         �                 � � �           u m     ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                   ��$     ����X� 06`	     �     N   N   n�     06`	N                  2         �                 � � �           u m     ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                   ��$     ����X� 06`	     �     N   N   n�     06`	N                  2         �                 � � �           u m     ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                   ��$     ����X� 06`	     �     N   N   n�     06`	N                  2         �                 � � �           u m     ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                   ��$     ����X� 06`	     �     N   N   n�     06`	N                  2         �                 � � �           u m     ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                   ��$     ����X� 06`	     �     N   N   n�     06`	N                  2         �                 � � �           u m     ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                   ��$     ����X� 06`	     �     N   N   n�     06`	N                  2         �                 � � �           u m     ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                   ��$     ����X� 06`	     �     N   N   n�     06`	N                  2         �                 � � �           u m     ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                   ��$     ����X� 06`	     �     N   N   n�     06`	N                  2         �                 � � �           u m     ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                   ��$     ����X� 06`	     �     N   N   n�     06`	N                  2         �                 � � �           u m     ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                   ��$     ����X� 06`	     �     N   N   n�     06`	N                  2         �                 � � �           u m     ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                   ��$     ����X� 06`	     �     N   N   n�     06`	N                  2         �                 � � �           u m     ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                   ��$     ����X� 06`	     �     N   N   n�     06`	N                  2         �                 � � �           u m     ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                   ��$     ����X� 06`	     �     N   N   n�     06`	N                  2         �                 � � �           u m     ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                   ��$     ����X� 06`	     �     N   N   n�     06`	N                  2         �                 � � �           u m     ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                   ��$     ����X� 06`	     �     N   N   n�     06`	N                  2         �                 � � �           u m     ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                   ��$     ����X� 06`	     �     N   N   n�     06`	N                  2         �                 � � �           u m     ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                   ��$     ����X� 06`	     �     N   N   n�     06`	N                  2         �                 � � �           u m     ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                   ��$     ����X� 06`	     �     N   N   n�     06`	N                  2         �                 � � �           u m     ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                   ��$     ����X� 06`	     �     N   N   n�     06`	N                  2         �                 � � �           u m     ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                   ��$     ����X� 06`	     �     N   N   n�     06`	N                  2         �                 � � �           u m     ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                   ��$     ����X� 06`	     �     N   N   n�     06`	N                  2         �                 � � �           u m     ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                   ��$     ����X� 06`	     �     N   N   n�     06`	N                  2         �                 � � �           u m     ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                   ��$     ����X� 06`	     �     N   N   n�     06`	N                  2         �                 � � �           u m     ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                               �� 	 CTitleBox                                                      �	                  @�         �  @                  ���                                                  �  @  B�     <   �  <     ��                                                        B�     |   �  |     ��                                                        B�     �   �  �     ��    � <                                                 B�     �   �  �     ��                                                        K� h      t  4     ��                                                      h      t  4   h      t  4   [title]                                       K� �   H   �  x     ��                                                      �   H   �  x   �   H   �  x   [description]                                       K� P   �   X  �     ��                                                      P   �   X  �   P   �   X  �   [id]                                       K� �   �   �  �     ��                                                      �   �   �  �   �   �   �  �   
[designer]                                       K�      ]   1    ��        	                                                   ]   1       ]   1  Date :       �	  4  �
  �                  K� p     x  4   	 ��        
                                              p     x  4  p     x  4  [date]                                       K�       U   1    
 ��                                                            U   1         U   1   Title :       �	  4  �
  �                  K�    L   �   q     ��                                                         L   �   q      L   �   q   Description :       �	  �  �  �                  K�    �   8   �     ��                                                         �   8   �      �   8   �   ID :       �	  �  8
  J                  K�    �   �   �     ��                                                         �   �   �      �   �   �   
Designer :       �	  t  p  
                   ��������������          �     	title box     Miscellaneous      �?    9 
 ��  CParamSubBehavior    
 R�  ����        ��������R�  ����       ��������R�  ����       ��������R�  ����       ��������R�  ����       ��������R�  ����       ��������R�  ����       ��������R�  ����       ��������R�  ����       ��������R�  ����  	     ��������        9                                      ������   CParamSubModelType�� ����  
   ��  	 CParmDefn            title                ��            description                ��            id                ��            designer                ��            Date :                ��            date                ��            Title :                ��            Description :                ��            ID :                ��            
Designer :                            ����             `         �?�� 	 CGraphDoc�  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                                                                                            2         �                 � � �                   ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                         U1Q2Q1Q0In1                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                      1m  0                            100   100                                                           1m  0                            100   100                              1m  0                            100   100                              1m  0                            100   100                                                 
               1m  0                            100   100                            ��   CPartPackage     ��   CPackage@  DO14�14 pin small outline package                                                                                                                                                                                                                              ����   yz{|}~   ���� ��@  DO14�14 pin small outline package                                                                                                                                                                                                                              ����   �����   ���q� ��@  DO14�14 pin small outline package                                                                                                                                                                                                                              ����   ������   � ��   CMiniPartPin    ����JJ     INJ�      ��   ����CkCk     INCk�     ��   ����KK     INK�     ��   ����RR     INR�     ��   ����QQ     OUTQ�     ��   ����Q'Q'     OUTQ'�          ��   CPackagePin 10 RIN 
 BB.Rƃ 1 JIN  AJƃ 4 KIN  AKƃ 8 JIN  BB.Jƃ 11 KIN  BB.Kƃ 3 QOUT  AA.Qƃ 2 Q'OUT  AA.Q'ƃ 13 RIN  AA.Rƃ 5 QOUT  BB.Qƃ 6 Q'OUT  BB.Q'ƃ 9 CkIN 	 BB.Clkƃ 12 CkIN  AA.ClkJK Flip-Flop w/clear
Flip FlopsGenericC      74107 A74107DA1               DIP1474107D74107D��  CXSpiceBehavior       jkclkresetoutnout ��   CBehPin     j����    �  j����                         ��Ճ    k����   �  k����                         ��Ճ    clk����   �  clk����                         ��Ճ     set����   �  set����                         ��Ճ    reset����   �  reset����                         ��Ճ    out����   �  out����                        ��Ճ    nout����   �  nout����                        ��74107 (XSpice)74107 (XSpice)  8               �������Digital<   Generic               ����    * time value noutQ'jJkKresetRoutQclkCk CkclkJjKkQ'noutQoutRreset                                                     � ��    ����JJ     INJ�      ��   ����CkCk     INCk�     ��   ����KK     INK�     ��   ����RR     INR�     ��   ����QQ     OUTQ�     ��   ����Q'Q'     OUTQ'�          ������������JK Flip-Flop w/clear
Flip FlopsGenericC      74107 A74107DA1               DIP1474107D74107DӃ       jkclkresetoutnout Ճ     j����    �  j����                         ��Ճ    k����   �  k����                         ��Ճ    clk����   �  clk����                         ��Ճ     set����   �  set����                         ��Ճ    reset����   �  reset����                         ��Ճ    out����   �  out����                        ��Ճ    nout����   �  nout����                        ��74107 (XSpice)74107 (XSpice)  8               �������Digital<   Generic               ����    * time value noutQ'jJkKresetRoutQclkCk CkclkJjKkQ'noutQoutRreset                                                     � ��    ����JJ     INJ�      ��   ����CkCk     INCk�     ��   ����KK     INK�     ��   ����RR     INR�     ��   ����QQ     OUTQ�     ��   ����Q'Q'     OUTQ'�      Z   ƃ 10 RPassive 
 BB.Rƃ 1 JIN  AJƃ 4 KIN  AKƃ 8 JPAS  BB.Jƃ 11 KPAS  BB.Kƃ 3 QOUT  AA.Qƃ 2 Q'OUT  AA.Q'ƃ 13 RIN  AA.Rƃ 5 QPassive  BB.Qƃ 6 Q'PAS  BB.Q'ƃ 9 CkPassive 	 BB.Clkƃ 12 CkIN  AA.ClkJK Flip-Flop w/clear
Flip FlopsGenericC      74107 A74107DA2                DIP1474107D74107DӃ       jkclkresetoutnout Ճ     j����    �  j����                         ��Ճ    k����   �  k����                         ��Ճ    clk����   �  clk����                         ��Ճ     set����   �  set����                         ��Ճ    reset����   �  reset����                         ��Ճ    out����   �  out����                        ��Ճ    nout����   �  nout����                        ��74107 (XSpice)74107 (XSpice)  8               �� Digital<   Generic               ����    * time value noutQ'jJkKresetRoutQclkCk CkclkJjKkQ'noutQoutRreset                                                     � ��    ����inIn     PAS1A�      ��   ����outY     PAS1Y�         ƃ 1 inPAS  A1Aƃ 2 outPAS  A1Yƃ 3 inPAS  B2Aƃ 4 outPAS  B2Yƃ 5 inPAS  C3Aƃ 6 outPAS  C3Yƃ 7  GND  COMGNDƃ 8 outPAS  D4Yƃ 9 inPAS 	 D4Aƃ 10 outPAS 
 E5Yƃ 11 inPAS  E5Aƃ 12 outPAS  F6Yƃ 13 inPAS  F6Aƃ 14  VCC  COMVCCdigital one-bit-wide inverterGatesGeneric=      7404 A7404DA3                                DIP147404D7404DӃ       inout Ճ     in����    �  in����                         ��Ճ    out����   �  out����                        ��7404 LS Inverter7404 LS Inverter  8               Digital<   Generic               ����    * time value inInoutY IninYout                        ��    ����AA     INA�      ClockClock                  ��    ����portport       ��������Output_PortOutput_Port                  ��    ����portport       ��������Output_PortOutput_Port                  ��    ����portport       ��������Output_PortOutput_Port                  ��    ����AA     INA      InputInput                  ��    ����aA     INaE      ��   ����bB     INbD     ��   ����cC     INcF     ��   ����yY     OUTyC     74ALS11A74ALS11A                                                                                 