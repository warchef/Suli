    � B2SPICE zzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzz    ��   TInPort        _   @         _   @                 Input��  CIntPin    ��  CWire      �         ��  CPart       �      p      �      p              74LS192D �   �    
 �      �	       �   �  p      �   �  p              74LS32D�    �    �        �       _   @         _   @                 Input ��  CExtPin    ��  CVertex          ��  CSegment    �2          �   �(   �      �   �,   �       �    �    `	          	                             �    �3      �    �     �   `  �   !                                        @  �   A     �  `          Up/Down     ��   CPin                    ��                                                       �   @   A��  TEllipse �   8   �   H                  ����
[negative]               ���                    �   8   �   H   �   8   �   H   �� 
 TRectangle t       �   @                   ����A                                      t       �   @   '� t   @   �   `                   ����A                                      t   @   �   `   ��  TLine �   @   �   @     ��                                                        '�         �   `                   ����                                                 �   `   *� t       t   `     
 ��                                                      ��  TPolygon                    ��                                                       ��  TPoint�   \        0��   P        0��   P        0��   D        0��   D        0��   P        0��   P    H�    .�                    ��                                                       0��   $        0��   0        0��   0        0��   <        0��   <        0��   0        0��   0    (�    ��  
 TTextField �       �   8    	 ��        	                                               �       �   8   �       �   8   	[A.nbits]      <       ����            �      "Arial                �       �   8   @�    (      M     ��        
                                                 (      M      (      M   [value]       �  �  $  n     (   l   P   @� ���������   #     ��                                                       ���������   #   ���������   #   	[refname]       �  Q  z  �  ���������       $ ,   +   ) 8   B / A C (   & -      input_general     Miscellaneous      �?      ��   TInPortModel       A ��  	 TModelPin Q  A����        A����                         ��             0��    ��������             0��    ��������             0��    ��������             0��    ��������             0��    ��������             0��    �������� d   :�0�yE>10e-9��    �������� d   :�0�yE>10e-9��    ��������                            ����  ����:�0�yE>10e-9��d         ����  ����:�0�yE>10e-9��d   �      E   �����        d   :�0�yE>10e-9��    �������� d   :�0�yE>10e-9��    ��������1 Bit Inport1 Bit Inport                 G Digital<   Generic   Up/DownUp/Down           ����  ��    �������� ����  ��    �������� ����  ��    �������� ����  ��    �������� ����  ��    �������� ����  ��    �������� ����  ��    ��������          ����            In ��   CPartPin    ����AA      INAA����    Digital Instruments Generic                         `   `              `   �  �              `   �             �  `   `          �      23  �        �         �  �        �  �              74LS04DJ �   �    �   M   �
       �   �  p      �   �  p              74LS32D�    �    �    Q    ��   TClock       �   �  �      �   �  �              ClockR �    �   �  �   �   V �   @  �   W �   �0   @  �   �   Z �/    	  �   [ �   �1    	  �   �   ^ �   `	  �   _    	        ]     \     �   \ �4    	  @   a �
   b �   `	  @   c    
                         Y     X                        �     A     �  �          Clock     #�                   ��                                                       �   `   A'�     @   �   �                  ����                                             @   �   �   *� �   `   �   `     ��                                                        *� `   @   `   �     ��                                                        *� p   h   x   h     ��    ����                                                *� x   T   x   h     ��    �                                                *� x   T   �   T     ��    ����                                                *� �   T   �   h     ��    �                                                  *� �   h   �   h     ��                                                        *� �   P   �   p      ��        	                                                @�    P   Z   u    
 ��        
                                                  P   m   u      P   m   u   [period]         p  (       P   P   t   @� �   `   �   �    	 ��                                                      �   `   �   �   �   `   �   �   ns       �  �  0  6  �   `   �   x   @�     �����        ��                                                           �����          �����      	[devname]        ����������������    �����      @�        X   @     ��                                                              X   @          X   @   	[refname]       �  �  �  h         �   <    n   m   l   k   j p   o q r i   h   g   e     f      Clock     Miscellaneous      �?      ��   TClockModel     ��  CValue '  ���ư>1000n      ��������u� �  ���Ơ>500n     �������� A F� �  A����        A����                          ��      x��    ��������      x��    ��������      x��    ��������      x��    ��������      x��    ��������      x��    �������� d   :�0�yE>10e-9��    �������� d   :�0�yE>10e-9��    ��������                             ����  ����:�0�yE>10e-9��d         ����  ����:�0�yE>10e-9��d   �     Q t   �����        d   :�0�yE>10e-9��    �������� d   :�0�yE>10e-9��    ��������ClockClock   �          x Digital InstrumentsO   Generic   ClockClock           ����  ��    �������� ����  ��    �������� ����  ��    �������� ����  ��    �������� ����  ��    �������� ����  ��    �������� ����  ��    ��������  lə    ����Generic            U H�    ����AA      INAA����    Digital InstrumentsDigital Clock inputGeneric                                                                             XH�                                   22 �   Q    22 P  x F�   B����       B����                          ��             0��    ��������             0��    ��������             0��    ��������             0��    ��������             0��    ��������             0��    �������� d   :�0�yE>10e-9��    �������� d   :�0�yE>10e-9��    ��������                             ����  ����:�0�yE>10e-9��d         ����  ����:�0�yE>10e-9��d   �     Q ��   TOr       ABY F�   A����        A����                          ��      x��    ��������      x��    ��������      x��    ��������      x��    ��������      x��    ��������      x��    �������� d   :�0�yE>10e-9��    �������� d   :�0�yE>10e-9��    ��������                             ����  ����:�0�yE>10e-9��d         ����  ����:�0�yE>10e-9��d   �      }   �����     ��   d   :�0�yE>10e-9��    �������� d   :�0�yE>10e-9��    ��������{ F�   Y����       Y����                         �� �   g5_P�W>22ns��    ��������      x��    �������� �   ��C֔N>14ns��    �������� �   g5_P�W>22ns��    ��������      x��    �������� �   ��C֔N>14ns��    �������� d   :�0�yE>10e-9��    �������� d   :�0�yE>10e-9��    ��������                            ����  ����:�0�yE>10e-9��d         ����  ����:�0�yE>10e-9��d   �      }   �����        d   :�0�yE>10e-9��    �������� d   :�0�yE>10e-9��    ��������32/4 LS 2-Inp. Or32/4 LS 2-Inp. Or  M 6i            ~ {  Digital<   Analog Devices   A2A2           ���� x��    �������� ���� x��    �������� @ �h㈵��>20u��    �������� ���-C��6:�-.4m��    �������� ���-C��6:�-.4m��    ��������  ������Mb�?8m��    ��������  Zb����Mbp?4m��    ��������   d     ����LS      �����     ��   d   :�0�yE>10e-9��    �������� d   :�0�yE>10e-9��    ��������F�   A����        A����                          ��      x��    ��������      x��    ��������      x��    ��������      x��    ��������      x��    ��������      x��    �������� d   :�0�yE>10e-9��    �������� d   :�0�yE>10e-9��    ��������                             ����  ����:�0�yE>10e-9��d         ����  ����:�0�yE>10e-9��d   �     Q |�       ABY � F�   B����       B����                          ��             0��    ��������             0��    ��������             0��    ��������             0��    ��������             0��    ��������             0��    �������� d   :�0�yE>10e-9��    �������� d   :�0�yE>10e-9��    ��������                             ����  ����:�0�yE>10e-9��d         ����  ����:�0�yE>10e-9��d   �     M �   �����     ��   d   :�0�yE>10e-9��    �������� d   :�0�yE>10e-9��    ��������F�   Y����       Y����                         �� �   g5_P�W>22ns��    ��������      x��    �������� �   ��C֔N>14ns��    �������� �   g5_P�W>22ns��    ��������      x��    �������� �   ��C֔N>14ns��    �������� d   :�0�yE>10e-9��    �������� d   :�0�yE>10e-9��    ��������                            ����  ����:�0�yE>10e-9��d         ����  ����:�0�yE>10e-9��d   �     �    �   �   	 28 �   �   O 28  F� �  Down����       Down����                          ��      x��    ��������      x��    ��������      x��    ��������      x��    ��������      x��    ��������      x��    �������� d   :�0�yE>10e-9��    �������� d   :�0�yE>10e-9��    ��������                            ����  ����:�0�yE>10e-9��d         ����  ����:�0�yE>10e-9��d   �     � ��   T74192       ClrUpDownLoadABCDCOBOQAQBQCQD F� �  Clr����        Clr����                          ��      x��    ��������      x��    ��������      x��    ��������      x��    ��������      x��    ��������      x��    �������� d   :�0�yE>10e-9��    �������� d   :�0�yE>10e-9��    ��������                             ����  ����:�0�yE>10e-9��d         ����  ����:�0�yE>10e-9��d   �      �   �����     ��   d   :�0�yE>10e-9��    �������� d   :�0�yE>10e-9��    ��������F� �  Up����       Up����                          ��      x��    ��������      x��    ��������      x��    ��������      x��    ��������      x��    ��������      x��    �������� d   :�0�yE>10e-9��    �������� d   :�0�yE>10e-9��    ��������                            ����  ����:�0�yE>10e-9��d         ����  ����:�0�yE>10e-9��d   �      �   �����     ��   d   :�0�yE>10e-9��    �������� d   :�0�yE>10e-9��    ��������� F� �  Load����       Load����                          ��      x��    ��������      x��    ��������      x��    ��������      x��    ��������      x��    ��������      x��    �������� d   :�0�yE>10e-9��    �������� d   :�0�yE>10e-9��    ��������                            ����  ����:�0�yE>10e-9��d         ����  ����:�0�yE>10e-9��d   �     �    �    �    �       _   @         _   @                 Input� �    �      �   �   � �7    
  �   � �   � �   @      �                               @  �   A     �  �          Load     #�                    ��                                                       �   @   A%� �   8   �   H                  ����
[negative]               ���                    �   8   �   H   �   8   �   H   '� t       �   @                   ����A                                      t       �   @   '� t   @   �   `                   ����A                                      t   @   �   `   *� �   @   �   @     ��                                                        '�         �   `                   ����                                                 �   `   *� t       t   `     
 ��                                                      .�                    ��                                                       0��   \        0��   P        0��   P        0��   D        0��   D        0��   P        0��   P    |�    .�                    ��                                                       0��   $        0��   0        0��   0        0��   <        0��   <        0��   0        0��   0    �|�    @� �       �   8    	 ��        	                                               �       �   8   �       �   8   	[A.nbits]      <       ����            �      "Arial                �       �   8   @�    (      M     ��        
                                                 (      M      (      M   [value]       �  8  $  �     (   l   P   @� ��������H   #     ��                                                       ��������H   #   ��������H   #   	[refname]       �  �  �  Q  ���������       � �   �   � �   � � � � �   � �      input_general     Miscellaneous      �?      D�       A F� Q  A����        A����                         ��             0��    ��������             0��    ��������             0��    ��������             0��    ��������             0��    ��������             0��    �������� d   :�0�yE>10e-9��    �������� d   :�0�yE>10e-9��    ��������                            ����  ����:�0�yE>10e-9��d         ����  ����:�0�yE>10e-9��d   �     � �   �����        d   :�0�yE>10e-9��    �������� d   :�0�yE>10e-9��    ��������1 Bit Inport1 Bit Inport   �            � Digital<   Generic   LoadLoad           ����  ��    �������� ����  ��    �������� ����  ��    �������� ����  ��    �������� ����  ��    �������� ����  ��    �������� ����  ��    ��������          ����            In H�    ����AA      INAA�<      Digital Instruments Generic                         `   `              `   �  �              `   �             �  `   `          �      11 �   �   	 11  � �  11�   �����     ��   d   :�0�yE>10e-9��    �������� d   :�0�yE>10e-9��    ��������F� �  A����       A����                          ��      x��    ��������      x��    ��������      x��    ��������      x��    ��������      x��    ��������      x��    �������� d   :�0�yE>10e-9��    �������� d   :�0�yE>10e-9��    ��������                             ����  ����:�0�yE>10e-9��d         ����  ����:�0�yE>10e-9��d   �     �    �    �    �       _   @         _   @                 Input� �   �    � �   �    ��   TBus       _      �      _      �              Splitter 1-to-4�    �    � 3  � �   �    �   �    � 5 � �   �   � 5  �   �   	 5  F� ����A:2����       A����                                        0��    ��������             0��    ��������             0��    ��������             0��    ��������             0��    ��������             0��    �������� d   :�0�yE>10e-9��    �������� d   :�0�yE>10e-9��    ��������                             ����  ����:�0�yE>10e-9��d         ����  ����:�0�yE>10e-9��d   �     � D�       A F� ����A:0����        A����                                         0��    ��������             0��    ��������             0��    ��������             0��    ��������             0��    ��������             0��    �������� d   :�0�yE>10e-9��    �������� d   :�0�yE>10e-9��    ��������                             ����  ����:�0�yE>10e-9��d         ����  ����:�0�yE>10e-9��d   �     � �   �����         d   :�0�yE>10e-9��    �������� d   :�0�yE>10e-9��    ��������F� ����A:1����       A����                                        0��    ��������             0��    ��������             0��    ��������             0��    ��������             0��    ��������             0��    �������� d   :�0�yE>10e-9��    �������� d   :�0�yE>10e-9��    ��������                             ����  ����:�0�yE>10e-9��d         ����  ����:�0�yE>10e-9��d   �     � �   �����        d   :�0�yE>10e-9��    �������� d   :�0�yE>10e-9��    ��������� F� ����A:3����       A����                                        0��    ��������             0��    ��������             0��    ��������             0��    ��������             0��    ��������             0��    �������� d   :�0�yE>10e-9��    �������� d   :�0�yE>10e-9��    ��������                             ����  ����:�0�yE>10e-9��d         ����  ����:�0�yE>10e-9��d   �     �    �   �    � 6 �   �    � 6  �   �   � 6  �   �   	 6  � F� �  D����       D����                          ��      x��    ��������      x��    ��������      x��    ��������      x��    ��������      x��    ��������      x��    �������� d   :�0�yE>10e-9��    �������� d   :�0�yE>10e-9��    ��������                             ����  ����:�0�yE>10e-9��d         ����  ����:�0�yE>10e-9��d   �     � �   �����     ��   d   :�0�yE>10e-9��    �������� d   :�0�yE>10e-9��    �������� 6�   �����         d   :�0�yE>10e-9��    �������� d   :�0�yE>10e-9��    ��������1 Bit Inport1 Bit Inport                 � � � � Digital<   Generic   ValueValue           ����  ��    �������� ����  ��    �������� ����  ��    �������� ����  ��    �������� ����  ��    �������� ����  ��    �������� ����  ��    ��������          ����            �����        d   :�0�yE>10e-9��    �������� d   :�0�yE>10e-9��    ��������F� �  C����       C����                          ��      x��    ��������      x��    ��������      x��    ��������      x��    ��������      x��    ��������      x��    �������� d   :�0�yE>10e-9��    �������� d   :�0�yE>10e-9��    ��������                             ����  ����:�0�yE>10e-9��d         ����  ����:�0�yE>10e-9��d   �     � �   �����     ��   d   :�0�yE>10e-9��    �������� d   :�0�yE>10e-9��    �������� 5   � 5  � �   �   � 3  �   �   � 4  � � �    �    `  �   �   �       
   �            �                       `   in    �   �   �  �   �   � �   @  �   �                        `   out1   �   �   �  �   �   � �   @      �                        �   out2   �   �&   �  @   �   � �	   @  �   �                           out3   �   �'   �  �   �   � �
   @  �   �                        �  out4    `             U2     #�                   ��                                                               in#�                   ��                                                      `       out1#�                   ��                                                      `   @   out2#�                   ��                                                      `   `   out3#�                    ��                                                      `   �   out4*� @       `         ��                                                      *� @   @   `   @     ��                                                      *� @   `   `   `     ��                                                      *� @   �   `   �     ��                                                      *�         @        	 ��        	                                              *�     @   @   @    
 ��        
                                              *�     `   @   `     ��                                                      *�     �   @   �     ��                                                      *�             �     ��                                                      @� D   d   N   }     ��                                                       D   d   N   }   D   d   N   }   [out4.bits]      <       ����            �      Times New Roman,  L  L  �  D   d   l   |   @� D   D   N   ]     ��                                                       D   D   N   ]   D   D   N   ]   [out3.bits]      <       ����            �      Times New Roman,  �  L  P  D   D   l   \   @� D   $   N   =     ��                                                       D   $   N   =   D   $   N   =   [out2.bits]      <       ����            �      Times New Roman,  �  L  �  D   $   h   <   @� D      N        ��                                                       D      N      D      N      [out1.bits]      <       ����            �      Times New Roman,  ,  L  �  D      l      @� ����            ��                                                       ����          ����          
[in.nbits]      <       ����            �      Times New RomanT     t  �  ����    (       �   �   � � � � � � � � � � �   � � �   � � �      busout4     Miscellaneous      �?      ��  	 CBehavior          bus 4bus 4  �             MiscellaneousY   Generic   U2U2            U  Wire Combiners & splitters Generic                                                                                                                                                                    4  � �   �   	 4  � F� �  B����       B����                          ��      x��    ��������      x��    ��������      x��    ��������      x��    ��������      x��    ��������      x��    �������� d   :�0�yE>10e-9��    �������� d   :�0�yE>10e-9��    ��������                             ����  ����:�0�yE>10e-9��d         ����  ����:�0�yE>10e-9��d   �     � �   �����     ��   d   :�0�yE>10e-9��    �������� d   :�0�yE>10e-9��    �������� 4   � 4 � � �    �    @  �   AQ   �  `	          Value     #�                    ��                                                       �   @   A%� �   8   �   H                  ����
[negative]               ���                    �   8   �   H   �   8   �   H   '� t       �   @                   ����A                                      t       �   @   '� t   @   �   `                   ����A                                      t   @   �   `   *� �   @   �   @     ��                                                        '�         �   `                   ����                                                 �   `   *� t       t   `     
 ��                                                      .�                    ��                                                       0��   \        0��   P        0��   P        0��   D        0��   D        0��   P        0��   P    H�    .�                    ��                                                       0��   $        0��   0        0��   0        0��   <        0��   <        0��   0        0��   0    (�    @� �       �   9    	 ��        	                                               �       �   9   �       �   9   	[A.nbits]      <       ����            �      "Arial�  �	  �  $
  �       �   8   @�    (      M     ��        
                                                 (      M      (      M   [value]       �  �	  $  n
     (   l   P   @� ��������S   #     ��                                                       ��������S   #   ��������S   #   	[refname]       �  Q	  �  �	  ���������       �        �   �      input_general     Miscellaneous      �?      �   In H�    ����AA       A         H�   ����AA      A <      H�   ����AA      A        H�   ����AA      A        Digital Instruments Generic                 �?       `   `              `   �  �              `   �              �  `   `          �      3 � � �   �   	 3  � �  3�   �����     ��   d   :�0�yE>10e-9��    �������� d   :�0�yE>10e-9��    ��������� � � F� �  CO����       CO����                         �� �   �A:��Y>24ns��    ��������      x��    �������� �   h�+e�SS>18ns��    ��������   �?Y��[>26ns��    ��������      x��    �������� �   �C���@R>17ns��    �������� d   :�0�yE>10e-9��    �������� d   :�0�yE>10e-9��    ��������                           ����  ����:�0�yE>10e-9��d         ����  ����:�0�yE>10e-9��d   �     �	    �    	 	 16 �      	 ��   TOutPort       _   @         _   @                 Output_Port�    �   �  @   �#   �   `  �   $ 	      #     	              �   port     �  �          Carry     #�                   ��                                                           @   port'�         �   `                   ����                                                 �   `   *�     @       @      ��                                                        %�    8       H                  ����
[negative]               ���                       8       H      8       H   @� (   ,   :   Q     ��                                                      (   ,   :   Q   (   ,   :   Q   [value]       8    p  �  (   ,   �   T   @�     $       <     ��                                                           $       <       $       <   [port.nbits]      <       ����            �      "Arial                    $       <   @�     ����r         ��                                                           ����r           ����r       	[refname]          h          �����       (  &)*+,'     Output_Port     Miscellaneous      �?      ��   TOutPortModel       port F� ����port����        port����                                         0��    ��������             0��    ��������             0��    ��������             0��    ��������             0��    ��������             0��    �������� d   :�0�yE>10e-9��    �������� d   :�0�yE>10e-9��    ��������                             ����  ����:�0�yE>10e-9��d         ����  ����:�0�yE>10e-9��d   �     .  �����     ��   d   :�0�yE>10e-9��    �������� d   :�0�yE>10e-9��    ��������Output_PortOutput_Port   �            /Digital<   Generic   CarryCarry           ����  ��    �������� ����  ��    �������� ����  ��    �������� ����  ��    �������� ����  ��    �������� ����  ��    �������� ����  ��    ��������  X{�    ����       ����  Out H�    ����portport       A   (     Digital Instruments Generic                                                                                                             16  /	 16�   �����        d   :�0�yE>10e-9��    �������� d   :�0�yE>10e-9��    ��������F� �  BO����	       BO����                         �� �   �A:��Y>24ns��    ��������      x��    �������� �   ,i�)+P>15ns��    �������� �   �A:��Y>24ns��    ��������      x��    �������� �   ��&�.Q>16ns��    �������� d   :�0�yE>10e-9��    �������� d   :�0�yE>10e-9��    ��������                           ����  ����:�0�yE>10e-9��d         ����  ����:�0�yE>10e-9��d   �     �
    �	   2	 
 	 17 �    2  
  �       _   @         _   @                 Output_Port4�    �   �  �   �$   �   `  @   8 
     	 7     
              �   port     �  �          Borrow     #�                   ��                                                           @   port'�         �   `                   ����                                                 �   `   *�     @       @      ��    ����                                                %�    8       H                  ����
[negative]               ���                       8       H      8       H   @� (   ,   :   Q     ��                                                      (   ,   :   Q   (   ,   :   Q   [value]       8  D  p  �  (   ,   �   T   @�     $       <     ��                                                           $       <       $       <   [port.nbits]      <       ����            �      "Arial                    $       <   @�     �����         ��                                                           �����           �����       	[refname]          �  `  H      �����       <  :=>?@;     Output_Port     Miscellaneous      �?      -�       port F� ����port����        port����                                         0��    ��������             0��    ��������             0��    ��������             0��    ��������             0��    ��������             0��    �������� d   :�0�yE>10e-9��    �������� d   :�0�yE>10e-9��    ��������                             ����  ����:�0�yE>10e-9��d         ����  ����:�0�yE>10e-9��d   �     2A  �����     ��   d   :�0�yE>10e-9��    �������� d   :�0�yE>10e-9��    ��������Output_PortOutput_Port   �            BDigital<   Generic   BorrowBorrow           ����  ��    �������� ����  ��    �������� ����  ��    �������� ����  ��    �������� ����  ��    �������� ����  ��    �������� ����  ��    ��������          ����       ����  Out H�    ����portport       A ��      Digital Instruments Generic                                                                           ����                                17  B1
 17�   �����        d   :�0�yE>10e-9��    �������� d   :�0�yE>10e-9��    ��������F� �  QA����
       QA����                         �� �  +�|�;i>47ns��    ��������      x��    ��������   �?Y��[>26ns��    �������� �  :�0�ye>40ns��    ��������      x��    �������� �   ����ba[>25.5ns��    �������� d   :�0�yE>10e-9��    �������� d   :�0�yE>10e-9��    ��������                            ����  ����:�0�yE>10e-9��d         ����  ����:�0�yE>10e-9��d   �     �    �
   E
  	 18 �   E  ��       _      �      _      �              Combiner 4-to-1�    E   H18  �   �    �   K  	 19 �   K  H19  J�   K    �       _   @         _   @                 Output_Port�    E   O18 N�   �    �   R  	 20 �   R  H20  �   R   H20  Q F� ����port:2����       port����                                        0��    ��������             0��    ��������             0��    ��������             0��    ��������             0��    ��������             0��    �������� d   :�0�yE>10e-9��    �������� d   :�0�yE>10e-9��    ��������                             ����  ����:�0�yE>10e-9��d         ����  ����:�0�yE>10e-9��d   �     R-�       port F� ����port:0����        port����                                         0��    ��������             0��    ��������             0��    ��������             0��    ��������             0��    ��������             0��    �������� d   :�0�yE>10e-9��    �������� d   :�0�yE>10e-9��    ��������                             ����  ����:�0�yE>10e-9��d         ����  ����:�0�yE>10e-9��d   �     EW  �����     ��   d   :�0�yE>10e-9��    �������� d   :�0�yE>10e-9��    ��������F� ����port:1����       port����                                        0��    ��������             0��    ��������             0��    ��������             0��    ��������             0��    ��������             0��    �������� d   :�0�yE>10e-9��    �������� d   :�0�yE>10e-9��    ��������                             ����  ����:�0�yE>10e-9��d         ����  ����:�0�yE>10e-9��d   �     KW  �����     ��   d   :�0�yE>10e-9��    �������� d   :�0�yE>10e-9��    ��������VF� ����port:3����       port����                                        0��    ��������             0��    ��������             0��    ��������             0��    ��������             0��    ��������             0��    �������� d   :�0�yE>10e-9��    �������� d   :�0�yE>10e-9��    ��������                             ����  ����:�0�yE>10e-9��d         ����  ����:�0�yE>10e-9��d   �     �    �   [  	 21 �   [  H21  �   [   H21  �   [   O21  ZF� �  QD����       QD����                         �� �  +�|�;i>47ns��    ��������      x��    ��������   �?Y��[>26ns��    �������� �  :�0�ye>40ns��    ��������      x��    �������� �   ����ba[>25.5ns��    �������� d   :�0�yE>10e-9��    �������� d   :�0�yE>10e-9��    ��������                            ����  ����:�0�yE>10e-9��d         ����  ����:�0�yE>10e-9��d   �     [�   �����        d   :�0�yE>10e-9��    �������� d   :�0�yE>10e-9��    �������� 21W  �����     ��   d   :�0�yE>10e-9��    �������� d   :�0�yE>10e-9��    ��������Output_PortOutput_Port   �            XYVZDigital<   Generic   OutputOutput           ����  ��    �������� ����  ��    �������� ����  ��    �������� ����  ��    �������� ����  ��    �������� ����  ��    �������� ����  ��    ��������          ����       ����  �����     ��   d   :�0�yE>10e-9��    �������� d   :�0�yE>10e-9��    ��������F� �  QC����       QC����                         �� �  +�|�;i>47ns��    ��������      x��    ��������   �?Y��[>26ns��    �������� �  :�0�ye>40ns��    ��������      x��    �������� �   ����ba[>25.5ns��    �������� d   :�0�yE>10e-9��    �������� d   :�0�yE>10e-9��    ��������                            ����  ����:�0�yE>10e-9��d         ����  ����:�0�yE>10e-9��d   �     R�   �����         d   :�0�yE>10e-9��    �������� d   :�0�yE>10e-9��    �������� 20   O20 _�    �   �      �"   �!   @  �   d           c                      �   port     �  `          Output     #�                   ��                                                           @   port'�         �   `                   ����                                                 �   `   *�     @       @      ��    ����                                                %�    8       H                  ����
[negative]               ���                       8       H      8       H   @� (   ,   :   Q     ��                                                      (   ,   :   Q   (   ,   :   Q   [value]       8  �  p  z  (   ,   �   T   @�     $   
   =     ��                                                           $   
   =       $   
   =   [port.nbits]      <       ����            �      "Arial�  �  �  0      $       <   @�     �����         ��                                                           �����           �����       	[refname]          H  X  �      �����       h  fijklg     Output_Port     Miscellaneous      �?      W  Out H�    ����portport       A  & -    H�   ����portport      A n Q   H�   ����portport      A �      H�   ����portport      A ��    Digital Instruments Generic                                                                           ����                                19  YF� �  QB����       QB����                         �� �  +�|�;i>47ns��    ��������      x��    ��������   �?Y��[>26ns��    �������� �  :�0�ye>40ns��    ��������      x��    �������� �   ����ba[>25.5ns��    �������� d   :�0�yE>10e-9��    �������� d   :�0�yE>10e-9��    ��������                            ����  ����:�0�yE>10e-9��d         ����  ����:�0�yE>10e-9��d   �     K�   �����         d   :�0�yE>10e-9��    �������� d   :�0�yE>10e-9��    �������� 19   H19  U^GMT]�    e      `   out    �   �"      �   �   �   `  �   u      
 t                 `   in1   �   �#          �   �   `      y       x                 �   in2   �   �$      �   �    �   `  �   }       |                    in3   �   �%      �   �!   �   `  �   �       �                 �  in4       `          U3     #�                    ��                                                       `       out#�                   ��                                                              in1#�                   ��                                                          @   in2#�                   ��                                                          `   in3#�                   ��                                                          �   in4*�                   ��                                                      *�     @       @     ��                                                      *�     `       `     ��                                                      *�     �       �     ��                                                      *�         `        	 ��        	                                              *�     @   @   @    
 ��        
                                              *�     `   @   `     ��                                                      *�     �   @   �     ��                                                      *� @       @   �     ��                                                      @�    d      }     ��                                                          d      }      d      }   
[in4.bits]      <       ����            �      Times New Roman8  �  X  �     d   0   |   @�    D      ]     ��                                                          D      ]      D      ]   
[in3.bits]      <       ����            �      Times New Roman8  ,  X  �     D   0   \   @�    $      =     ��                                                          $      =      $      =   
[in2.bits]      <       ����            �      Times New Roman8  �  X  0     $   ,   <   @�               ��                                                                               
[in1.bits]      <       ����            �      Times New Roman8  l  X  �        0      @� H      R        ��                                                       H      R      H      R      [out.nbits]      <       ����            �      Times New Roman�  l    �  H      t       ��  �  ���������������  �     busin4     Miscellaneous      �?      ��          bus 4bus 4  �             MiscellaneousY   Generic   U3U3            U  Wire Combiners & splitters Generic                                                                                                                                                                    18  IP XD 18�   �����         d   :�0�yE>10e-9��    �������� d   :�0�yE>10e-9��    ��������qa`192 LS Up/Down Counter192 LS Up/Down Counter  b 6i            � � � � � � � � 1Dqa`Digital<   Generic   A1A1           ���� x��    �������� ���� x��    �������� @ �h㈵��>20u��    �������� ���-C��6:�-.4m��    �������� ���,C��6:�-400u��    ��������  ������Mb�?8m��    �������� �+S��~j�t�?19m��    ��������          ����LS     2   :�0�y5>5n��    �������� ����    ��~A32meg��    �������� �   :�0�yU>20n��    �������� �   �C���@R>17n��    ��������  �����     ��   d   :�0�yE>10e-9��    �������� d   :�0�yE>10e-9��    ���������  28�   �����        d   :�0�yE>10e-9��    �������� d   :�0�yE>10e-9��    ��������32/4 LS 2-Inp. Or32/4 LS 2-Inp. Or  M 6i            � � � Digital<   Analog Devices   A3A3           ���� x��    �������� ���� x��    �������� @ �h㈵��>20u��    �������� ���-C��6:�-.4m��    �������� ���-C��6:�-.4m��    ��������  ������Mb�?8m��    ��������  Zb����Mbp?4m��    ��������          ����LS      �����     ��   d   :�0�yE>10e-9��    �������� d   :�0�yE>10e-9��    �������� 22   O 22 N � �    d           aȇ��   �   `	      �   �6    	      �   �5    	  �   �   �   @  �   �       �    �    �    �    �       
          �  b   �   �   @  �   �   ��   @  @   �              
      �  �  y    `	             A3     #�                   ��                                                           `   a#�                   ��                                                          �   b#�                    ��                                                      �   �   y��   TArc    0   �   �    	                                                              0   �   �      0   �   �   D   �   �   �           *�     P   D   P     ��                                                        ��    P   �   �                                                                  P   �   �      P   �   �   �   �   D   P           *�     �   D   �     ��                                                        *� �   �   �   �     ��                                                        *�     `   ,   `     ��                                                        *�     �   ,   �     ��        	                                                ��    P   0   �    
           
                                                   P   0   �      P   0   �   $   �   $   P           @�     (   B   P     ��                                                           (   B   P       (   B   P   	[refname]       `	  �  (
  8      (   t   L   @�        �   (     ��                                                              �   (          �   (   	[devname]        ����������������       �   (    �  ����  �  ����  �  �  �     OR 2    	OR 2 IEEEMiscellaneous      �?    M  �   A H�    ����aA      INA1A�>      H�   ����bB      INA1B�>     H�   ����yY      OUTA1Y�>     H�    ����aA      INB1A�>      H�   ����bB      INB1B�>     H�   ����yY      OUTB1Y����   H�    ����aA      INC1A�>      H�   ����bB      INC1B�>     H�   ����yY      OUTC1Y����   H�    ����aA      IND1A����    H�   ����bB      IND1B����   H�   ����yY      OUTD1Y����   Gatesdigital n-input OR gateGenericDO14             27 L  � F� 8  Y����       Y����                         �� �   ,i�)+P>15ns��    ��������      x��    �������� d   :�0�yE>10ns��    �������� �   ,i�)+P>15ns��    ��������      x��    �������� Z   h�+e�SC>9ns��    �������� d   :�0�yE>10e-9��    �������� d   :�0�yE>10e-9��    ��������                           ����  ����:�0�yE>10e-9��d         ����  ����:�0�yE>10e-9��d   �     M ��   TAnd       InY F� 7  In����        In����                          ��      x��    ��������      x��    ��������      x��    ��������      x��    ��������      x��    ��������      x��    �������� d   :�0�yE>10e-9��    �������� d   :�0�yE>10e-9��    ��������                             ����  ����:�0�yE>10e-9��d         ����  ����:�0�yE>10e-9��d   �      �  �����     ��   d   :�0�yE>10e-9��    �������� d   :�0�yE>10e-9��    ���������04/6 LS Inverter04/6 LS Inverter =               ��Digital<   Generic   A4A4           ���� x��    �������� ���� x��    �������� @ �h㈵��>20u��    �������� ���-C��6:�-.4m��    �������� ���-C��6:�-.4m��    ��������  ������Mb�?8m��    ��������  6nb2U0*�c?2.4m��    ��������          ����LS      �����         d   :�0�yE>10e-9��    �������� d   :�0�yE>10e-9��    �������� 27  K 27 �    "        �  in    �   �  �  �  out    `             A4     #�                   ��                                                           �   in#�                   ��                                                      �   �   out%� l   t   �   �                   ���                                          l   t   �   �   l   t   �   �   *� �   �   �   �     ��    ����                                                *�     �   ,   �     ��    ����                                                .� ����    ����      ��                                                         0�,   \    h��0�,   �    *a�L0�l   �       0�,   \            @� ����   �   0     ��                                                       ����   �   0   ����   �   0   	[devname]        ��������������������   �   0   @� ����0   >   X     ��                                                       ����0   >   X   ����0   >   X   	[refname]       T  �    P  ����0   �   T   	 �  �������     Inverter    Inverter IEEEMiscellaneous      �?    =  �  A H�    ����inIn      INA1AInpu    H�   ����outY      OUTA1Y      H�    ����inIn      INB1A       H�   ����outY      OUTB1Y      H�    ����inIn      INC1Azzzz    H�   ����outY      OUTC1Y       H�    ����inIn      IND1A  E    H�   ����outY      OUTD1Y1 B   H�    ����inIn      INE1A����    H�   ����outY      OUTE1Y  ��   H�    ����inIn      INF1AAA�    H�   ����outY      OUTF1Y       Gatesdigital one-bit-wide inverterGenericDO14              23  G ~ � 23    23 z  �               a    �   `       �  b   �   �-   @  `   �   ��+   `  `   ��   ��.   `  �   �	   ��   @  �   �           �                   	      �  �  y    `	  �          A2     #�                   ��                                                           `   a#�                   ��                                                          �   b#�                    ��                                                      �   �   y��    0   �   �    	                                                              0   �   �      0   �   �   D   �   �   �           *�     P   D   P     ��                                                        ��    P   �   �                                                                  P   �   �      P   �   �   �   �   D   P           *�     �   D   �     ��                                                        *� �   �   �   �     ��                                                        *�     `   ,   `     ��                                                        *�     �   ,   �     ��        	                                                ��    P   0   �    
           
                                                   P   0   �      P   0   �   $   �   $   P           @�     (   B   P     ��                                                           (   B   P       (   B   P   	[refname]       `	  X  (
  �      (   t   L   @�        �   (     ��                                                              �   (          �   (   	[devname]        ����������������       �   (    �  ����  �  ����  �  �  �     OR 2    	OR 2 IEEEMiscellaneous      �?    M  }   A H�    ����aA      INA1A 0��    H�   ����bB      INA1B       H�   ����yY      OUTA1Y       H�    ����aA      INB1A�      H�   ����bB      INB1B     H�   ����yY      OUTB1Y       H�    ����aA      INC1A       H�   ����bB      INC1B      H�   ����yY      OUTC1Y       H�    ����aA      IND1A       H�   ����bB      IND1B     H�   ����yY      OUTD1Y     Gatesdigital n-input OR gateGenericDO14              25  �   25  	 25 � � � � � 3FLS\�    �   @      �    �)   �      �   �*   �  @   �   �      @                                                    �  Clr    �   �      �  Up   �   �      �  Down   �   �       `  Load   �   �          A   �   �       �  B   �   �       �  C   �   �       @  D   �   %     �  CO   �	   9 	    �  BO	   �
   v 
       QA
   �   z     �  QB   �   ~     �  QC   �   �     @  QD    @  �          A1    A #�                   ��                                                           �   Clr#�                   ��                                                          �   Up#�                   ��                                                          �   Down#�                   ��                                                             Load#�                   ��                                                          `  A#�                   ��                                                          �  B#�                   ��                                                          �  C#�                   ��                                                          �  D#�                  	 ��                                                      `  �   CO#�                  
 ��        	                                              `  �   BO#�                   ��        
                                              `  `  QA#�                   ��                                                      `  �  QB#�                   ��                                                      `  �  QC#�                   ��                                                      `  �  QD'� @   P     �                 ����                                         @   P     �  *�     �   @   �     ��                                                        *�     �   @   �     ��                                                        *�     �   @   �     ��                                                        *�    �   4  �    . ��                                                        *�    �      �    / ��                                                        *�     �           3 ��                                                        *�        @       2 ��                                                        *�     �   @   �    1 ��                                                        *�     �       �    0 ��                                                        *� @   p     p   6 ��                                                        *� @   �     �   7 ��                                                        *� @   �     �   8 ��                                                        *� �   �   �   �    = ��                                                        *� �   �   �   �    > ��                                                        *�        @        ��                                                        *�     `  @   `    ��    (O�                                                *�     �  @   �    ��                                                        *�     �  @   �    ��                                                         *�     �  @   �    ��        !                                                *�    �   `  �     ��        "                                                *�    �   `  �     ��        #                                                *�    `  `  `    ��        $                                                *�    �  `  �    ��        %                                                *�    �  `  �    ��        &                                                *�    �  `  �    ��        '                                                *� @   �   L   �    & ��        (                                                *� L   �   @   �    ' ��        )                                                *� L   �   @   �    ( ��        *                                                *� @   �   L   �    ) ��        +                                                *� ,     ,       * ��        ,                                                *� ,     @       + ��        -                                                *�    �   4  �    , ��       .                                                *�    �      �    - ��    ���/                                                .� ����������������   ��        0                                                 0�P   P  0 �ݙ0�P   @  0 �ݙ0�@   @  0 �ݙ0�@   @   0 �ݙ0�   @   0 �ݙ0�   @  0 �ݙ0�  @  0 �w�0�  P  0 �ݙ    @� H   p   �   �     ��        1                                              H   p   �   �   H   p   �   �   ct=0         �  �  �  H   p   �   �   @� T   �   y   �     ��        2                                              T   �   y   �   T   �   y   �   2+       <  P  �  �  T   �   |   �   @� T   �   q   �      ��        3                                              T   �   q   �   T   �   q   �   1-       <    �  �  T   �   |   �   @� H     j   5   ! ��        4                                              H     j   5  H     j   5  c3         �  �  f  H     �   0  @� H   P  m   u   " ��        5                                              H   P  m   u  H   P  m   u  3d         �  �  &  H   P  t   p  @� h   @   �   e    # ��        6                                              h   @   �   e   h   @   �   e   	ctrdIv 10       x  `  �  �  h   @     `   @� H   �   m   �    4 ��        7                                              H   �   m   �   H   �   m   �   g1         �  �  F  H   �   p   �   @� �   �     �    $ ��        8                                              �   �     �   �   �     �   1ct=9       �  P  p  �  �   �      �   @� �   �     �    % ��        9                                              �   �     �   �   �     �   2ct=0       �    p  �  �   �      �   @� H   �   m      5 ��        :                                              H   �   m     H   �   m     g2         p  �    H   �   p     @� �   L  �   q   9 ��        ;                                              �   L  �   q  �   L  �   q  [1]       ,  �  �    �   L  �   l  @� �   l  �   �   : ��        <                                              �   l  �   �  �   l  �   �  [2]       ,  �  �  z  �   l  �   �  @� �   �  �   �   ; ��        =                                              �   �  �   �  �   �  �   �  [4]       ,  D  �  �  �   �  �   �  @� �   �  �   �   < ��        >                                              �   �  �   �  �   �  �   �  [8]       ,  �  �  :  �   �  �   �  @� @      j   <    ? ��        ?                                               @      j   <   @      j   <   	[refname]          �  �  |  @      �   8   @� @   �����       @ ��        @                                               @   �����      @   �����      	[devname]        ����������������@   �����      c D   !"#$%123456789:MNOPQRTU;                <=>?@AVBSCWXYZ    [\                                  &'+  *  )  ,-.(      /0�     74192 Up/Down Counter     Miscellaneous      �?    b  �   A H�    ����ClrClr      INACLR�<      H�   ����UpUp      INAUP�<     H�   ����DownDown      INADOWN�<     H�   ����LoadLoad      INA~LOAD�<     H�   ����AA      INAA�<     H�   ����BB      INAB�<     H�   ����CC      INAC�<     H�   ����DD      INAD�<     H�   ����COCO      OUTA~CO�<     H�	   ����BOBO      OUTA~BO�<  	   H�
   ����QAQA      OUTAQA�<  
   H�   ����QBQB      OUTAQB�<     H�   ����QCQC      OUTAQC       H�   ����QDQD      OUTAQD       Counters(synchronous 4-bit up/down decade counterGenericDO16              8  F� Q  A����        A����                         ��             0��    ��������             0��    ��������             0��    ��������             0��    ��������             0��    ��������             0��    �������� d   :�0�yE>10e-9��    �������� d   :�0�yE>10e-9��    ��������                            ����  ����:�0�yE>10e-9��d         ����  ����:�0�yE>10e-9��d   �      D�       A k1 Bit Inport1 Bit Inport   �            kDigital<   Generic   ResetReset           ����  ��    �������� ����  ��    �������� ����  ��    �������� ����  ��    �������� ����  ��    �������� ����  ��    �������� ����  ��    ��������  ��    ����             �����         d   :�0�yE>10e-9��    �������� d   :�0�yE>10e-9��    ���������   8  �� 8 �       @  �   A     �  �          Reset     #�                    ��                                                       �   @   A%� �   8   �   H                  ����
[negative]               ���                    �   8   �   H   �   8   �   H   '� t       �   @                   ����A                                      t       �   @   '� t   @   �   `                   ����A                                      t   @   �   `   *� �   @   �   @     ��                                                       '�         �   `                   ����                                                 �   `   *� t       t   `     
 ��    ՛�w                                              .�                    ��                                                       0��   \        0��   P        0��   P        0��   D        0��   D        0��   P        0��   P    p��    .�                    ��                                                       0��   $        0��   0        0��   0        0��   <        0��   <        0��   0        0��   0    0��    @� �       �   8    	 ��        	                                               �       �   8   �       �   8   	[A.nbits]      <       ����            �      "Arial                �       �   8   @�    (      M     ��        
                                                 (      M      (      M   [value]       �  �  $  �     (   l   P   @� ��������X   #     ��                                                       ��������X   #   ��������X   #   	[refname]       �  q  �    ���������       ns  r  q}  �u��p  ot,�    input_general     Miscellaneous      �?      l  In H�    ����AA      INAA�      Digital Instruments Generic                         `   `              `   �  �              `   �             �  `   `          �       � � 	 !5OT  O K � H     � � � � �  � 2EKR[Q M % % %    W ���c a Y _   ! [ ] ��� �� � �� � � � uy}�d$8: 8 :   � � �� � � � � %9vz~�� #7cV X ` d ��" �� � � etx|�� �  � ��\ Z ^    b ���                  
 u�@ ����        ��������u�             0     ��������u� ����      @5     ��������u�  ʚ;�������?.1     ��������u�@ ����       ��������u� ����       ��������u� ����       ��������u� ����       ��������u� ���� true
     ��������u� ����  false     ��������               
                  u� ����        ��������u� ����       ��������u�  ����       ��������u�@ ����       ��������u�@ ����       ��������               
                  u� ����        ��������u� ����       ��������u�@ ����       ��������u�  ����       ��������u� ����       ��������u� ����       ��������u� ����       ��������u� ����       ��������u� ����       ��������u� ����       ��������u� ����       ��������               
                 u� ����dec     ��������u� ����     @�@1k     ��������u� ����    ��.A1meg     ��������u� ����       20     ��������u� ���� true     ��������u� ���� true     ��������u� ���� true	     ��������u� ����  false
     ��������               
                 u�  ����        ��������u�  ����       ��������u�  ����       ��������u� ����dec     ��������u� ����       ��������u� ����       ��������u� ����  	     ��������u� ����  
     ��������               
                  	 u� ����        ��������u� ����       ��������u� ����       ��������u� ����       ��������u� ����       ��������u� ����       ��������u� ����       ��������u� ����       ��������u� ����       ��������               
                 u� ����        ��������u� ����       ��������u� ����       ��������u� ����dec     ��������u� ����       ��������               
                     u�             0      ��������u� ��� ����MbP?1m     ��������u� �� �h㈵��>10u     ��������u� '  ���ư>1u     ��������u� ���� true     ��������u� ����  false     ��������u� ���� true     ��������u� ����  false     ��������               
                 u� ����     @�@1K      ��������u�  ����       ��������u�  ����       ��������u�  ����       ��������               
         ��              u�  ����        ��������              
                  u�  ����        ��������              
                                  
                 u�@ ����        ��������u�@ ����       ��������u� ����       ��������u� ����       ��������u� ����       ��������u� ����       ��������u� ����       ��������u� ����       ��������u� ����       ��������u� ���� true	     ��������u� ����  false
     ��������u� ���� true     ��������u� ����  false     ��������               
                 u� ����       5      ��������u� ����       5     ��������u� ����       5     ��������u� ����       5     ��������u� ����       ��������u� ����  	     ��������u� ����  
     ��������u� ����       ��������u� ����       ��������u� ����       ��������u� ���� true     ��������u�@ ����       ��������u�@ ����       ��������u� ����       ��������u� ����       ��������u� ����       ��������u� ����dec     ��������u� ����       ��������u� ����       ��������u� ����       ��������u� ���� true     ��������u� ���� true     ��������u� ���� true     ��������u� ����  false     ��������u� ���� true     ��������u� ����  false      ��������u� ���� true!     ��������u� ����  false"     ��������               
                        u� ����       5      ��������u� ����       5     ��������u� ����       5     ��������u� ����       5     ��������u� ����       ��������u� ����  	     ��������u� ����  
     ��������u� ����       ��������u� ����       ��������u� ����       ��������u� ���� true     ��������u�@ ����       ��������u�@ ����       ��������u� ����       ��������u� ����       ��������u� ����       ��������u� ����dec     ��������u� ����       ��������u� ����       ��������u� ����       ��������u� ���� true     ��������u� ���� true     ��������u� ���� true     ��������u� ����  false     ��������u� ���� true     ��������u� ����  false      ��������u� ���� true!     ��������u� ����  false"     ��������               
                 u� ����       5      ��������u� ����       5     ��������u� ����       5     ��������u� ����       5     ��������u� ����       ��������u� ����  	     ��������u� ����  
     ��������u� ����       ��������u� ����       ��������u� ����       ��������u� ���� true     ��������u�@ ����       ��������u�@ ����       ��������u� ����       ��������u� ����       ��������u� ����       ��������u� ����dec     ��������u� ����       ��������u� ����       ��������u� ����       ��������u� ���� true     ��������u� ���� true     ��������u� ���� true     ��������u� ����  false     ��������u� ���� true     ��������u� ����  false      ��������u� ���� true!     ��������u� ����  false"     ��������               
                 u� ����       5      ��������u� ����       5     ��������u� ����       5     ��������u� ����       5     ��������u� ����       ��������u� ����  	     ��������u� ����  
     ��������u� ����       ��������u� ����       ��������u� ����       ��������u� ���� true     ��������u�@ ����       ��������u�@ ����       ��������u� ����       ��������u� ����       ��������u� ����       ��������u� ����dec     ��������u� ����       ��������u� ����       ��������u� ����       ��������u� ���� true     ��������u� ���� true     ��������u� ���� true     ��������u� ����  false     ��������u� ���� true     ��������u� ����  false      ��������u� ���� true!     ��������u� ����  false"     ��������               
                 u�@ ����        ��������u�@ ����       ��������u� ����       ��������u� ����       ��������u� ����       ��������u� ����       ��������u� ����       ��������u� ����       ��������u� ����decade     ��������u� ���� true     ��������u� ���� true     ��������u� ���� true     ��������u� ����  false     ��������               
                 u� ����        ��������u� ����       ��������u�@ ����       ��������u�  ����       ��������u� ����       ��������u� ����       ��������u� ����       ��������u� ����       ��������u� ����       ��������u� ����       ��������u� ����       ��������               
                        u� ����dec     ��������u� ����     @�@1k     ��������u� ����    ��.A1meg     ��������u� ����       20     ��������u� ����        0     ��������u� ����        0     ��������u� ���� true	     ��������u� ���� true
     ��������u� ����      I@50     ��������u� ���� true     ��������u� ����  false     ��������               
                          / u� ���� x'     ��������u�     �-���q=1E-12     ��������u� @B -C��6?1E-4     ��������u� ���� x     ��������u� ���� x     ��������u� ���� x     ��������u� ���� x     ��������u� ���� x     ��������u� ���� x     ��������u� ���� x	     ��������u� ���� x!     ��������u� ����    �  500
     ��������u� ���� x     ��������u� ����    �  500     ��������u� ���� x$     ��������u� ���� x$     ��������u� ���� x%     ��������u� ���� x"     ��������u�  ���� x*     ��������u� ���� x     ��������u� ���� x     ��������u� ���� x     ��������u� ���� x&     ��������u� ���� x     ��������u� ���� x     ��������u� ���� x     ��������u� ���� x+     ��������u� ���� x,     ��������u� ���� x-     ��������u� ���� xg     ��������u� ���� xf     ��������u� ���� xd     ��������u� ���� xe     ��������u� ���� xh     ��������u� ���� xj     ��������u� ���� xi     ��������u� ���� xk     ��������u� ����    e��A1Gl     ��������u�             0�     ��������u� ����      @5�     ��������u� ����      @2.5�     ��������u� ����      �?.5�     ��������u� ����      @4.5�     ��������u� 
   ��&�.>1n�     ��������u� 
   ��&�.>1n�     ��������u� 
   ��&�.>1n�     ��������u� 
   ��&�.>1n�     ��������                                  Ariald        ��=i�px�  �=i,� ��/i    ��=i�px�  �=i,� ��/i ��  COpAnal                         
                        ����                                   ��=i�px�  �=i,� ��/i    ��=i�px�  �=i,� ��/i ��  CDCsweep       
 ����������               
                      ����                                   ��=i�px�  �=i,� ��/i    ��=i�px�  �=i,� ��/i ��  CACsweep        ��������               
                      ����                                  ��=i�px�  �=i,� ��/i    ��=i�px�  �=i,� ��/i �� 
 CTranSweep        ��������               
                      ����                                   ��=i�px�  �=i,� ��/i    ��=i�px�  �=i,� ��/i ��  CACdisto        �����               
                          ����                                  ��=i�px�  �=i,� ��/i    ��=i�px�  �=i,� ��/i ��        u� ����        ��������u� ����       ��������u� ����       ��������u� ����dec     ��������u� ����       ��������               
                          ����                                  ��=i�px�  �=i,� ��/i    ��=i�px�  �=i,� ��/i ��        u� ����        ��������u� ����       ��������u� ����       ��������u� ����dec     ��������u� ����       ��������               
                          ����                                  ��=i�px�  �=i,� ��/i    ��=i�px�  �=i,� ��/i ��        u� ����        ��������u� ����       ��������u� ����       ��������u� ����dec     ��������u� ����       ��������               
                          ����                                  ��=i�px�  �=i,� ��/i    ��=i�px�  �=i,� ��/i ��        u� ����        ��������u� ����       ��������u� ����       ��������u� ����dec     ��������u� ����       ��������               
                          ����           � �                    ��=i�px�  �=i,� ��/i    ��=i�px�  �=i,� ��/i ��        u� ����        ��������u� ����       ��������u� ����       ��������u� ����dec     ��������u� ����       ��������               
                      	    ����                                  ��=i�px�  �=i,� ��/i    ��=i�px�  �=i,� ��/i ��  CACnoise        ��������               
                   
    ����                                  ��=i�px�  �=i,� ��/i    ��=i�px�  �=i,� ��/i ƃ                        
                        ����                                  ��=i�px�  �=i,� ��/i    ��=i�px�  �=i,� ��/i ��  CFourier        ����               
         ��                  ����                                   ��=i�px�  �=i,� ��/i    ��=i�px�  �=i,� ��/i ��  CACpz        	 ���������               
                       ����                                   ��=i�px�  �=i,� ��/i    ��=i�px�  �=i,� ��/i ��  CDCtf         �����               
                       ����                                   ��=i�px�  �=i,� ��/i    ��=i�px�  �=i,� ��/i ��  CDCsens         �����������               
                       ����                                   ��=i�px�  �=i,� ��/i    ��=i�px�  �=i,� ��/i                 ����                                   ��=i�px�  �=i,� ��/i    ��=i�px�  �=i,� ��/i ��  CShow         �              
                       ����                                   ��=i�px�  �=i,� ��/i    ��=i�px�  �=i,� ��/i ��  CShowmod         �              
                       ����                                   ��=i�px�  �=i,� ��/i    ��=i�px�  �=i,� ��/i �� 
 CLinearize        u�  ����        ��������               
                      ����                                   ��=i�px�  �=i,� ��/i    ��=i�px�  �=i,� ��/i ��  CParamTranSweep        �������������               
                      ����                                   ��=i�px�  �=i,� ��/i    ��=i�px�  �=i,� ��/i �             ����                                   ��=i�px�  �=i,� ��/i    ��=i�px�  �=i,� ��/i ��  CParamACSweep        LMNOPQRSTUVWX               
                      ����                                  ��=i�px�  �=i,� ��/i    ��=i�px�  �=i,� ��/i ��  CMonteCarlo_op        ����������������������������               
                             ����                                   ��=i�px�  �=i,� ��/i    ��=i�px�  �=i,� ��/i ��  CMonteCarlo_dc        �������� 	
               
                      ����                                   ��=i�px�  �=i,� ��/i    ��=i�px�  �=i,� ��/i ��  CMonteCarlo_ac         !"#$%&'()*+,-./               
                      ����                                  ��=i�px�  �=i,� ��/i    ��=i�px�  �=i,� ��/i ��  CMonteCarlo_tran        0123456789:;<=>?@ABCDEFGHIJK               
                      ����                                   ��=i�px�  �=i,� ��/i    ��=i�px�  �=i,� ��/i ��  CACsens        YZ[\]^_`abc               
                             ����                                  ��=i�px�  �=i,� ��/i    ��=i�px�  �=i,� ��/i ��  CNetworkAnalysis        defghijklmn               
                      ����                                  ��=i�px�  �=i,� ��/i    ��=i�px�  �=i,� ��/i                 ����                                 >           ��   CDigSimResTemplate                           ��   TDigitalSignal            Reset    ���� ����                        �            Up/Down    ���� ����                        �            Value   ���� ����                        �            Load    ���� ����                        �            Carry    ���� ����                        �            Borrow    ���� ����                        �            Output   ���� ����                        �            Clock    ���� ����                                  ���       ����  ����:�0�yU>+20.00n���   ����                       Arial����                       Arial����                       Arial                                           ����  ���� ������       ����  ���� ������                 �               ����  �����       200������          0.000000e+000��    ��������      0.000000e+000��    ��������      0.000000e+000��    ��������   ����                       Arial����                       Arial����                       Arial����                       Arial                        �     �   �  �                     ����  ��    ��������                                                         A  DO16�16 pin small outline package                                                                                                                                                                                                                              ����   ��   CPackageAliasSuperPCBStandardSO16      �EagleBURR.LBRSO16-1      �Orcad SOG.050/16/WG.255/L.400      �Pads SO16NB      �	UltiboardL7IC.l55$SO16      �Eaglesmd-ipc.lbrSO16             A                                                                                    @  DO14�14 pin small outline package                                                                                                                                                                                                                              ����   �SuperPCBStandardSO14      �EagleBURR.LBRSO14      �Orcad SOG.050/14/WG.244/L.350      �Pads SO14NB      �	UltiboardL7IC.l55$SO14      �Eagleburr-brown.lbrSO14             A        @  DO14�14 pin small outline package                                                                                                                                                                                                                              ����   ������        B        @  DO14�14 pin small outline package                                                                                                                                                                                                                              ����   �SuperPCBStandardSO14      �EagleBURR.LBRSO14      �Orcad SOG.050/14/WG.244/L.350      �Pads SO14NB      �	UltiboardL7IC.l55$SO14      �Eagleburr-brown.lbrSO14             A                        �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                   ط�     ����t� �w    <�     h   h   ��     �wh                  2         �                 � � �           k t     ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                   ط�     ����t� �w    <�     h   h   ��     �wh                  2         �                 � � �           k t     ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                   ط�     ����t� �w    <�     h   h   ��     �wh                  2         �                 � � �           k t     ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                   ط�     ����t� �w    <�     h   h   ��     �wh                  2         �                 � � �           k t     ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                   ط�     ����t� �w    <�     h   h   ��     �wh                  2         �                 � � �           k t     ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                   ط�     ����t� �w    <�     h   h   ��     �wh                  2         �                 � � �           k t     ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                   ط�     ����t� �w    <�     h   h   ��     �wh                  2         �                 � � �           k t     ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                   ط�     ����t� �w    <�     h   h   ��     �wh                  2         �                 � � �           k t     ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                   ط�     ����t� �w    <�     h   h   ��     �wh                  2         �                 � � �           k t     ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                   ط�     ����t� �w    <�     h   h   ��     �wh                  2         �                 � � �           k t     ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                   ط�     ����t� �w    <�     h   h   ��     �wh                  2         �                 � � �           k t     ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                   ط�     ����t� �w    <�     h   h   ��     �wh                  2         �                 � � �           k t     ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                   ط�     ����t� �w    <�     h   h   ��     �wh                  2         �                 � � �           k t     ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                   ط�     ����t� �w    <�     h   h   ��     �wh                  2         �                 � � �           k t     ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                   ط�     ����t� �w    <�     h   h   ��     �wh                  2         �                 � � �           k t     ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                   ط�     ����t� �w    <�     h   h   ��     �wh                  2         �                 � � �           k t     ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                   ط�     ����t� �w    <�     h   h   ��     �wh                  2         �                 � � �           k t     ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                   ط�     ����t� �w    <�     h   h   ��     �wh                  2         �                 � � �           k t     ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                   ط�     ����t� �w    <�     h   h   ��     �wh                  2         �                 � � �           k t     ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                   ط�     ����t� �w    <�     h   h   ��     �wh                  2         �                 � � �           k t     ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                   ط�     ����t� �w    <�     h   h   ��     �wh                  2         �                 � � �           k t     ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                   ط�     ����t� �w    <�     h   h   ��     �wh                  2         �                 � � �           k t     ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                   ط�     ����t� �w    <�     h   h   ��     �wh                  2         �                 � � �           k t     ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                   ط�     ����t� �w    <�     h   h   ��     �wh                  2         �                 � � �           k t     ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                   ط�     ����t� �w    <�     h   h   ��     �wh                  2         �                 � � �           k t     ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                   ط�     ����t� �w    <�     h   h   ��     �wh                  2         �                 � � �           k t     ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                   ط�     ����t� �w    <�     h   h   ��     �wh                  2         �                 � � �           k t     ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                   ط�     ����t� �w    <�     h   h   ��     �wh                  2         �                 � � �           k t     ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                   ط�     ����t� �w    <�     h   h   ��     �wh                  2         �                 � � �           k t     ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                   ط�     ����t� �w    <�     h   h   ��     �wh                  2         �                 � � �           k t     ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                               �� 	 CTitleBox                                                      �	                  '�         �  @                  ���                                                  �  @  *�     <   �  <     ��                                                        *�     |   �  |     ��                                                        *�     �   �  �     ��                                                        *�     �   �  �     ��                                                        @� h      t  4     ��                                                      h      t  4   h      t  4   [title]                                       @� �   H   �  x     ��                                                      �   H   �  x   �   H   �  x   [description]                                       @� P   �   X  �     ��                                                      P   �   X  �   P   �   X  �   [id]                                       @� �   �   �  �     ��                                                      �   �   �  �   �   �   �  �   
[designer]                                       @�      ]   1    ��        	                                                   ]   1       ]   1  Date :       �  4  �  �                  @� p     x  4   	 ��        
                                              p     x  4  p     x  4  [date]                                       @�       U   1    
 ��                                                            U   1         U   1   Title :       �  4  �  �                  @�    L   �   q     ��                                                         L   �   q      L   �   q   Description :       �  �  �   �                  @�    �   8   �     ��                                                         �   8   �      �   8   �   ID :       �  �  8  J                  @�    �   �   �     ��                                                         �   �   �      �   �   �   
Designer :       �  t  p   
                   	
               	title box     Miscellaneous      �?    9 
 ��  CParamSubBehavior    
 u�  ����        ��������u�  ����       ��������u�  ����       ��������u�  ����       ��������u�  ����       ��������u�  ����       ��������u�  ����       ��������u�  ����       ��������u�  ����       ��������u�  ����  	     ��������        9                                      ������   CParamSubModelType�� ����  
   ��  	 CParmDefn            title                %�            description                %�            id                %�            designer                %�            Date :                %�            date                %�            Title :                %�            Description :                %�            ID :                %�            
Designer :                            ����             `         �?�� 	 CGraphDoc�  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                                                                                            2         �                 � � �                   ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                         ResetUp/DownValueLoadCarryBorrowOutputClock                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                      1m  0                            100   100                                                           1m  0                            100   100                              1m  0                            100   100                              1m  0                            100   100                                                 
               1m  0                            100   100                            ��   CPartPackageࣣ ��   CPackageA  DO16�16 pin small outline package                                                                                                                                                                                                                              ����   ������   2�|�� 4�@  DO14�14 pin small outline package                                                                                                                                                                                                                              ����   ������   2��k� 4�@  DO14�14 pin small outline package                                                                                                                                                                                                                              ����          ��   CMiniPartPin    ����AA     INA  Q  InputInput                  :�    ����AA     INA  Q  InputInput                  :�    ����AA       ��������:�   ����AA      ��������:�   ����AA      ��������:�   ����AA      ��������InputInput                              :�    ����AA     INA  Q  InputInput               3 :�    ����ClrClr     INCLR�  �<  :�   ����UpUp     INUP�  �<  :�   ����DownDown     INDOWN 	  �<  :�   ����LoadLoad     IN~LOAD	  �<  :�   ����AA     INA	  �<  :�   ����BB     INB	  �<  :�   ����CC     INC	  �<  :�   ����DD     IND	  �<  :�   ����COCO     OUT~CO	  �<  :�	   ����BOBO     OUT~BO	  �<  :�
   ����QAQA     OUTQA	  �<  :�   ����QBQB     OUTQB		  �<  :�   ����QCQC     OUTQC
	  �<  :�   ����QDQD     OUTQD	  �<   	   ��   CPackagePin 14 Clr   ACLRP� 5 Up   AUPP� 4 Down   ADOWNP� 11 Load   A~LOADP� 15 A   AAP� 1 B   ABP� 10 C  
 ACP� 9 D  	 ADP� 12 CO   A~COP� 13 BO   A~BOP� 3 QA   AQAP� 2 QB   AQBP� 6 QC   AQCP� 7 QD   AQDP� 8  GND  COMGNDP� 16  VCC  COMVCC(synchronous 4-bit up/down decade counterCountersGenericF      74192 A74LS192DA1            DIP1674LS192D74LS192D��  CXSpiceBehavior       clrupdownloadabcdcoboqaqbqcqd ��   CBehPin �<  clr����    u  clr����                         ��c� �<  up����   u  up����                         ��c� �<  down����   u  down����                         ��c� �<  load����   u  load����                         ��c� �<  a����   u  a����                        ��c� �<  b����   u  b����                         ��c� �<  c����   u  c����                         ��c� �<  d����   u  d����                        ��c� �<  co����   u  co����                        ��c� �<  bo����	   u  bo����                        ��c� �<  qa����
   u  qa����                       ��c� �<  qb����   u  qb����                        ��c� �<  qc����   u  qc����                        ��c� �<  qd����   u  qd����                       ��74192 LS (XSpice)74192 LS (XSpice)  8 �            defghijklmnopqDigital<   Generic                       * time value qaQAdownDownqbQBclrClrqcQCqdQDloadLoadupUpaAcoCObBboBOcCdD DdDowndownQAqaQBqbQCqcLoadloadQDqdClrclrUpupCOcoBOboAaBbCc                                                                                                                        :�    ����portport       ��������Output_PortOutput_Port                  :�    ����portport       ��������Output_PortOutput_Port                  :�    ����portport       ��������:�   ����portport      ��������:�   ����portport      ��������:�   ����portport      ��������Output_PortOutput_Port                              :�    ����AA     INA�  �  ClockClock               6 :�    ����aA     IN1A.  �Q  :�   ����bB     IN1B/  �Q  :�   ����yY     OUT1Y0  �Q    O   P� 1 a   A1AP� 2 b   A1BP� 3 y   A1YP� 4 a   B2AP� 5 b   B2BP� 6 y   B2YP� 7  GND  COMGNDP� 8 y   C3YP� 9 a  	 C3AP� 10 b  
 C3BP� 11 y   D4YP� 12 a   D4AP� 13 b   D4BP� 14  VCC  COMVCCdigital n-input OR gateGatesGeneric=      7432 A74LS32DA2                       DIP1474LS32D74LS32Da�       aby c� �Q  a����    �  a����                        ��c� �Q  b����   �  b����                        ��c� �Q  y����   �  y����                        ��74LS32 2-input Or74LS32 2-input Or  8               ���Digital<   Generic                       * time value yYaAbB YyAaBb                             6 :�    ����aA     IN1A.  �Q  :�   ����bB     IN1B/  �Q  :�   ����yY     OUT1Y0  �Q    O   |}~����������digital n-input OR gateGatesGeneric=      7432 A74LS32DA2                       DIP1474LS32D74LS32D                               8 :�    ����inIn     IN1A�  �>  :�   ����outY     OUT1Y�  �>   K   P� 1 in   A1AP� 2 out   A1YP� 3 in   B2AP� 4 out   B2YP� 5 in   C3AP� 6 out   C3YP� 7  GND  COMGNDP� 8 out   D4YP� 9 in  	 D4AP� 10 out  
 E5YP� 11 in   E5AP� 12 out   F6YP� 13 in   F6AP� 14  VCC  COMVCCdigital one-bit-wide inverterGatesGeneric=      7404 A74LS04DA3                                DIP1474LS04D74LS04Da�       inout c� �>  in����    �  in����                         ��c� �>  out����   �  out����                        ��7404 LS Inverter7404 LS Inverter  8               ��Digital<   Generic                       * time value inInoutY IninYout                         Splitter 1-to-4Splitter 1-to-4                                                               Combiner 4-to-1Combiner 4-to-1                                                                                                     