    � B2SPICE zzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzz    ��  CPart          @  `        @  `              74LS109D��  CIntPin    ��  CWire      �         ��   TInPort       _   @         _   @                 Input ��  CExtPin    ��  CVertex&      �   ��  CSegment    �#   �  �   �    �   �                      �    �$      �   �    �                         �    �"   �  �   �'    �   �                     �2    �?   �  �    �3    �!   �       �4    �@   �  `                                                                          @  �   A     �              In2     ��   CPin                    ��                                                       �   @   A��  TEllipse �   8   �   H                  ����
[negative]               ���                    �   8   �   H   �   8   �   H   �� 
 TRectangle t       �   @                   ����A                                      t       �   @   %� t   @   �   `                   ����A                                      t   @   �   `   ��  TLine �   @   �   @     ��                                                        %�         �   `                   ����                                                 �   `   (� t       t   `     
 ��                                                      ��  TPolygon                    ��                                                       ��  TPoint�   \        .��   P        .��   P        .��   D        .��   D    ��  .��   P        .��   P    �ʁ    ,�                    ��                                                       .��   $        .��   0        .��   0    �Ut.��   <    tY.��   <     ���.��   0      9�.��   0    `�z    ��  
 TTextField �       �   8    	 ��        	                                               �       �   8   �       �   8   	[A.nbits]      <       ����            �      "Arial                �       �   8   >�    (      M     ��        
                                                 (      M      (      M   [value]       �   x         (   l   P   >� ��������+   #     ��                                                       ��������+   #   ��������+   #   	[refname]       �   �  B  �  ���������       " *   )   ' 6   @ - ? A &   $ +      input_general     Miscellaneous      �?      ��   TInPortModel       A ��  	 TModelPin Q  A����        A����                         ��             0��    ��������             0��    ��������             0��    ��������             0��    ��������             0��    ��������             0��    �������� d   :�0�yE>10e-9��    �������� d   :�0�yE>10e-9��    ��������                            ����  ����:�0�yE>10e-9��d         ����  ����:�0�yE>10e-9��d   �      C   �����        d   :�0�yE>10e-9��    �������� d   :�0�yE>10e-9��    ��������1 Bit Inport1 Bit Inport                 E Digital<   Generic   In2In2           ����  ��    �������� ����  ��    �������� ����  ��    �������� ����  ��    �������� ����  ��    �������� ����  ��    �������� ����  ��    ��������          ����            In ��   CPartPin    ����AA      INAA�      Digital Instruments Generic                         `   `              `   �  �              `   �   t�z       �  `   `          �      14 �         �         @  `        @  `              74LS109DH �   �    �   K    12 J �   K   I 12 �   K   �         @  `        @  `              74LS109D�         O 14 N �   �    �   R    3 �    R    ��   TClock       �   �  �      �   �  �              ClockT 
�    �   �  �
   �   X �    `  �
   Y �
   Z �   @  �
   �   �   @      �   ^ �	          _            ]     \     [ �	   \ �      �
   �   �          c �   d �   �      e                b     a �   b �7      �
   g �   �8          i �   j �
   `      k �   l �9   �      m                        h                             �   �   `      �   p �   �      q             o     Z                        �     A     �  �	          U1     !�                   ��                                                       �   `   A%�     @   �   �                  ����                                             @   �   �   (� �   `   �   `     ��                                                        (� `   @   `   �     ��                                                        (� p   h   x   h     ��                                                        (� x   T   x   h     ��                                                        (� x   T   �   T     ��                                                        (� �   T   �   h     ��                                                        (� �   h   �   h     ��                                                        (� �   P   �   p      ��        	                                                >�    P   Z   u    
 ��        
                                                  P   Z   u      P   Z   u   [period]         �
  �  F     P   P   t   >� �   `   �   �    	 ��                                                      �   `   �   �   �   `   �   �   ns       �  �
  0  v  �   `   �   x   >�     �����        ��                                                           �����          �����      	[devname]        ����������������    �����      >�        *   @     ��                                                              *   @          *   @   	[refname]       �  
  `  �
         �   <    |   {   z   y   x ~   }  � w   v   u   s     t      Clock     Miscellaneous      �?      ��   TClockModel     ��  CValue �  I�����z>100n      ���������� �  I�����j>50n     �������� A D� �  A����        A����                          ��      x��    ��������      x��    ��������      x��    ��������      x��    ��������      x��    ��������      x��    �������� d   :�0�yE>10e-9��    �������� d   :�0�yE>10e-9��    ��������                             ����  ����:�0�yE>10e-9��d         ����  ����:�0�yE>10e-9��d   �     R �   �����         d   :�0�yE>10e-9��    �������� d   :�0�yE>10e-9��    ��������ClockClock   l           � Digital InstrumentsO   Generic   U1U1           ����  ��    �������� ����  ��    �������� ����  ��    �������� ����  ��    �������� ����  ��    �������� ����  ��    �������� ����  ��    ��������          ����Generic             U F�    ����AA      INAA       Digital InstrumentsDigital Clock inputGeneric                                                                                                                   3 �   R   I 3 Q �   R   �         @  `        @  `              74LS109D�         � 14 �   �    �   �   O 16 � �    �    ��   TOutPort
       _   @         _   @                 Output_Port� 
�    �0   �  @   �(   � �/   �  �   � �   �   �  �   �        �     �/   � �   `  �   � �0   � �>   �  �   �                               
            �   port     �  �          Out3     !�                   ��                                                           @   port%�         �   `                   ����                                                 �   `   (�     @       @      ��    ����                                                #�    8       H                  ����
[negative]               ���                       8       H      8       H   >� (   ,   E   Q     ��                                                      (   ,   E   Q   (   ,   E   Q   [value]       �    P  �  (   ,   �   T   >�     $       <     ��                                                           $       <       $       <   [port.nbits]      <       ����            �      "Arial                    $       <   >�     ����j         ��                                                           ����j           ����j       	[refname]       �  h  �        �����       �   � � � � � �      Output_Port     Miscellaneous      �?      ��   TOutPortModel       port D� ����port����        port����                                         0��    ��������             0��    ��������             0��    ��������             0��    ��������             0��    ��������             0��    �������� d   :�0�yE>10e-9��    �������� d   :�0�yE>10e-9��    ��������                             ����  ����:�0�yE>10e-9��d         ����  ����:�0�yE>10e-9��d   �     � �   �����     ��   d   :�0�yE>10e-9��    �������� d   :�0�yE>10e-9��    ��������Output_PortOutput_Port                 � Digital<   Generic   Out3Out3           ����  ��    �������� ����  ��    �������� ����  ��    �������� ����  ��    �������� ����  ��    �������� ����  ��    �������� ����  ��    ��������          ����       ����  Out F�    ����portport       A �>      Digital Instruments Generic               SS                                                                                           16  � D� P  Q����       Q����                         �� �  :�0�ye>40ns��    ��������      x��    �������� �   I�����Z>25ns��    �������� �   I�����Z>25ns��    ��������      x��    �������� �   �?Y��K>13ns��    �������� d   :�0�yE>10e-9��    �������� d   :�0�yE>10e-9��    ��������                            ����  ����:�0�yE>10e-9��d         ����  ����:�0�yE>10e-9��d   �     � ��   TJKFF_general       SJClkKRQQ' D� K  S����        S����                          ��      x��    ��������      x��    ��������      x��    ��������      x��    ��������      x��    ��������      x��    �������� d   :�0�yE>10e-9��    �������� d   :�0�yE>10e-9��    ��������                            ����  ����:�0�yE>10e-9��d         ����  ����:�0�yE>10e-9��d   �      �   �����     ��   d   :�0�yE>10e-9��    �������� d   :�0�yE>10e-9��    ��������D� L  J����       J����                          ��      x��    ��������      x��    ��������      x��    ��������      x��    ��������      x��    ��������      x��    �������� d   :�0�yE>10e-9��    �������� d   :�0�yE>10e-9��    ��������                             ����  ����:�0�yE>10e-9��d         ����  ����:�0�yE>10e-9��d   �     K �   �����     ��   d   :�0�yE>10e-9��    �������� d   :�0�yE>10e-9��    ��������D� M  Clk����       Clk����                          ��      x��    ��������      x��    ��������      x��    ��������      x��    ��������      x��    ��������      x��    �������� d   :�0�yE>10e-9��    �������� d   :�0�yE>10e-9��    ��������                            ����  ����:�0�yE>10e-9��d         ����  ����:�0�yE>10e-9��d   �     R �   �����     ��   d   :�0�yE>10e-9��    �������� d   :�0�yE>10e-9��    ��������D� N  K����       K����                          ��      x��    ��������      x��    ��������      x��    ��������      x��    ��������      x��    ��������      x��    �������� d   :�0�yE>10e-9��    �������� d   :�0�yE>10e-9��    ��������                            ����  ����:�0�yE>10e-9��d         ����  ����:�0�yE>10e-9��d   �     �    �   �   I 7 �   �   O 7  D� Q  Q'����       Q'����                         �� �  :�0�ye>40ns��    ��������      x��    �������� �   I�����Z>25ns��    �������� �   I�����Z>25ns��    ��������      x��    �������� �   �?Y��K>13ns��    �������� d   :�0�yE>10e-9��    �������� d   :�0�yE>10e-9��    ��������                           ����  ����:�0�yE>10e-9��d         ����  ����:�0�yE>10e-9��d   �     � ��       SJClkKRQQ' D� K  S����        S����                          ��      x��    ��������      x��    ��������      x��    ��������      x��    ��������      x��    ��������      x��    �������� d   :�0�yE>10e-9��    �������� d   :�0�yE>10e-9��    ��������                            ����  ����:�0�yE>10e-9��d         ����  ����:�0�yE>10e-9��d   �      �   �����     ��   d   :�0�yE>10e-9��    �������� d   :�0�yE>10e-9��    ��������D� L  J����       J����                          ��      x��    ��������      x��    ��������      x��    ��������      x��    ��������      x��    ��������      x��    �������� d   :�0�yE>10e-9��    �������� d   :�0�yE>10e-9��    ��������                             ����  ����:�0�yE>10e-9��d         ����  ����:�0�yE>10e-9��d   �     K �   �����     ��   d   :�0�yE>10e-9��    �������� d   :�0�yE>10e-9��    ��������D� M  Clk����       Clk����                          ��      x��    ��������      x��    ��������      x��    ��������      x��    ��������      x��    ��������      x��    �������� d   :�0�yE>10e-9��    �������� d   :�0�yE>10e-9��    ��������                            ����  ����:�0�yE>10e-9��d         ����  ����:�0�yE>10e-9��d   �     R �   �����     ��   d   :�0�yE>10e-9��    �������� d   :�0�yE>10e-9��    ��������D� N  K����       K����                          ��      x��    ��������      x��    ��������      x��    ��������      x��    ��������      x��    ��������      x��    �������� d   :�0�yE>10e-9��    �������� d   :�0�yE>10e-9��    ��������                            ����  ����:�0�yE>10e-9��d         ����  ����:�0�yE>10e-9��d   �     �    �   �    13 �   �   I 13  D� Q  Q'����       Q'����                         �� �  :�0�ye>40ns��    ��������      x��    �������� �   I�����Z>25ns��    �������� �   I�����Z>25ns��    ��������      x��    �������� �   �?Y��K>13ns��    �������� d   :�0�yE>10e-9��    �������� d   :�0�yE>10e-9��    ��������                           ����  ����:�0�yE>10e-9��d         ����  ����:�0�yE>10e-9��d   �     � ��       SJClkKRQQ' D� K  S����        S����                          ��      x��    ��������      x��    ��������      x��    ��������      x��    ��������      x��    ��������      x��    �������� d   :�0�yE>10e-9��    �������� d   :�0�yE>10e-9��    ��������                            ����  ����:�0�yE>10e-9��d         ����  ����:�0�yE>10e-9��d   �      �   �����     ��   d   :�0�yE>10e-9��    �������� d   :�0�yE>10e-9��    ��������D� L  J����       J����                          ��      x��    ��������      x��    ��������      x��    ��������      x��    ��������      x��    ��������      x��    �������� d   :�0�yE>10e-9��    �������� d   :�0�yE>10e-9��    ��������                             ����  ����:�0�yE>10e-9��d         ����  ����:�0�yE>10e-9��d   �     �    �   �    4 �    �    �       _   @         _   @                 Input� �   �
    �  D� ����A:1����       A����                                        0��    ��������             0��    ��������             0��    ��������             0��    ��������             0��    ��������             0��    �������� d   :�0�yE>10e-9��    �������� d   :�0�yE>10e-9��    ��������                             ����  ����:�0�yE>10e-9��d         ����  ����:�0�yE>10e-9��d   �     � B�       A D� ����A:0����        A����                                         0��    ��������             0��    ��������             0��    ��������             0��    ��������             0��    ��������             0��    �������� d   :�0�yE>10e-9��    �������� d   :�0�yE>10e-9��    ��������                             ����  ����:�0�yE>10e-9��d         ����  ����:�0�yE>10e-9��d   �     � �   �����        d   :�0�yE>10e-9��    �������� d   :�0�yE>10e-9��    ��������� D� ����A:2����       A����                                        0��    ��������             0��    ��������             0��    ��������             0��    ��������             0��    ��������             0��    �������� d   :�0�yE>10e-9��    �������� d   :�0�yE>10e-9��    ��������                             ����  ����:�0�yE>10e-9��d         ����  ����:�0�yE>10e-9��d   �     �    �   �    � 9  �  9�   �����         d   :�0�yE>10e-9��    �������� d   :�0�yE>10e-9��    ��������D� ����A:3����       A����                                        0��    ��������             0��    ��������             0��    ��������             0��    ��������             0��    ��������             0��    �������� d   :�0�yE>10e-9��    �������� d   :�0�yE>10e-9��    ��������                             ����  ����:�0�yE>10e-9��d         ����  ����:�0�yE>10e-9��d   �     �    �   �    � 10  �  10�   �����         d   :�0�yE>10e-9��    �������� d   :�0�yE>10e-9��    ��������1 Bit Inport1 Bit Inport                 � � � � Digital<   Generic   SetSet           ����  ��    �������� ����  ��    �������� ����  ��    �������� ����  ��    �������� ����  ��    �������� ����  ��    �������� ����  ��    ��������          ����            �����         d   :�0�yE>10e-9��    �������� d   :�0�yE>10e-9��    ��������
 8  
 � 8 � � 
�    �          �*   � �      �   �   � �   �  �   �   
             � �   � �2      �   � �   � �   `  �   �   
               
           
           
            @  �   A     �   @          Set     !�                    ��                                                       �   @   A#� �   8   �   H                  ����
[negative]               ���                    �   8   �   H   �   8   �   H   %� t       �   @                   ����A                                      t       �   @   %� t   @   �   `                   ����A                                      t   @   �   `   (� �   @   �   @     ��                                                        %�         �   `                   ����                                                 �   `   (� t       t   `     
 ��                                                      ,�                    ��                                                       .��   \        .��   P        .��   P        .��   D        .��   D        .��   P        .��   P    �!w    ,�                    ��                                                       .��   $        .��   0        .��   0        .��   <        .��   <        .��   0        .��   0    p"w    >� �       �   9    	 ��        	                                               �       �   9   �       �   9   	[A.nbits]      <       ����            �      "Arial�  �  �    �       �   8   >�    (      M     ��        
                                                 (      M      (      M   [value]       �   �    N     (   l   P   >� ��������3   #     ��                                                       ��������3   #   ��������3   #   	[refname]       �   1  Z  �  ���������       � �   �   � �   � � � � �   � �      input_general     Miscellaneous      �?      �   In F�    ����AA       A ����    F�   ����AA      A �     F�   ����AA      A        F�   ����AA      A 0     Digital Instruments Generic                         `   `              `   �  �              `   �             �  `   `          �      4 �    �    �         �  �        �  �              74LS04D� �   �    �   �    5 �  D� N  K����       K����                          ��      x��    ��������      x��    ��������      x��    ��������      x��    ��������      x��    ��������      x��    �������� d   :�0�yE>10e-9��    �������� d   :�0�yE>10e-9��    ��������                            ����  ����:�0�yE>10e-9��d         ����  ����:�0�yE>10e-9��d   �     � �   �����     ��   d   :�0�yE>10e-9��    �������� d   :�0�yE>10e-9��    ��������D� 8  Y����       Y����                         �� �   ,i�)+P>15ns��    ��������      x��    �������� d   :�0�yE>10ns��    �������� �   ,i�)+P>15ns��    ��������      x��    �������� Z   h�+e�SC>9ns��    �������� d   :�0�yE>10e-9��    �������� d   :�0�yE>10e-9��    ��������                           ����  ����:�0�yE>10e-9��d         ����  ����:�0�yE>10e-9��d   �     � ��   TAnd       InY D� 7  In����        In����                          ��      x��    ��������      x��    ��������      x��    ��������      x��    ��������      x��    ��������      x��    �������� d   :�0�yE>10e-9��    �������� d   :�0�yE>10e-9��    ��������                             ����  ����:�0�yE>10e-9��d         ����  ����:�0�yE>10e-9��d   �     � �   �����     ��   d   :�0�yE>10e-9��    �������� d   :�0�yE>10e-9��    ��������� 04/6 LS Inverter04/6 LS Inverter =               � � Digital<   Generic   A4A4           ���� x��    �������� ���� x��    �������� @ �h㈵��>20u��    �������� ���-C��6:�-.4m��    �������� ���-C��6:�-.4m��    ��������  ������Mb�?8m��    ��������  6nb2U0*�c?2.4m��    ��������          ����LS      �����         d   :�0�yE>10e-9��    �������� d   :�0�yE>10e-9��    �������� 5  � 5 
�    �        �  in    
�   �1   @  �   �)   �   �  �                        �  �  out    `             A4     !�                   ��                                                           �   in!�                   ��                                                      �   �   out#� l   t   �   �                   ���                                          l   t   �   �   l   t   �   �   (� �   �   �   �     ��                                                        (�     �   ,   �     ��                                                        ,� ����    ����      ��                                                         .�,   \    ��v.�,   �        .�l   �    �Ut.�,   \            >� ����   �   0     ��                                                       ����   �   0   ����   �   0   	[devname]        ��������������������   �   0   >� ����0   >   X     ��                                                       ����0   >   X   ����0   >   X   	[refname]       T  �    0  ����0   �   T   	   	     Inverter    Inverter IEEEMiscellaneous      �?    =  �   A F�    ����inIn      INA1A�>      F�   ����outY      OUTA1Y�>     F�    ����inIn      INB1A d     F�   ����outY      OUTB1Y       F�    ����inIn      INC1A ���    F�   ����outY      OUTC1Y :�   F�    ����inIn      IND1A���:    F�   ����outY      OUTD1Y0e-9   F�    ����inIn      INE1A   7    F�   ����outY      OUTE1Y����   F�    ����inIn      INF1A�?8    F�   ����outY      OUTF1YinI   Gatesdigital one-bit-wide inverterGenericDO14              4  � � �  4�   �����     ��   d   :�0�yE>10e-9��    �������� d   :�0�yE>10e-9��    ��������D� M  Clk����       Clk����                          ��      x��    ��������      x��    ��������      x��    ��������      x��    ��������      x��    ��������      x��    �������� d   :�0�yE>10e-9��    �������� d   :�0�yE>10e-9��    ��������                            ����  ����:�0�yE>10e-9��d         ����  ����:�0�yE>10e-9��d   �     R �   �����     ��   d   :�0�yE>10e-9��    �������� d   :�0�yE>10e-9��    ��������� D� O  R����       R����                          ��      x��    ��������      x��    ��������      x��    ��������      x��    ��������      x��    ��������      x��    �������� d   :�0�yE>10e-9��    �������� d   :�0�yE>10e-9��    ��������                            ����  ����:�0�yE>10e-9��d         ����  ����:�0�yE>10e-9��d   �     �    �      11 �       �       _   @         _   @                 Input 
�    �%      �   �   #�'   �  �   �   �   �  @   &        %    $�   %�(      �   (�   �      @   *       )    �!   )�)   �  �   �   �   �  @   .       -    ,�    -�;   �  �   �+   �4   �  @   2       1    0                                           @  �   A     �              Reset     !�                    ��                                                       �   @   A#� �   8   �   H                  ����
[negative]               ���                    �   8   �   H   �   8   �   H   %� t       �   @                   ����A                                      t       �   @   %� t   @   �   `                   ����A                                      t   @   �   `   (� �   @   �   @     ��                                                        %�         �   `                   ����                                                 �   `   (� t       t   `     
 ��    ����                                              ,�                    ��                                                       .��   \        .��   P        .��   P     �� .��   D        .��   D        .��   P      ��.��   P    ��z    ,�                    ��                                                       .��   $        .��   0    (� t.��   0        .��   <        .��   <        .��   0       .��   0    `�z    >� �       �   8    	 ��        	                                               �       �   8   �       �   8   	[A.nbits]      <       ����            �      "Arial                �       �   8   >�    (      M     ��        
                                                 (      M      (      M   [value]       �   �    .     (   l   P   >� ��������X   #     ��                                                       ��������X   #   ��������X   #   	[refname]       �     �  �  ���������       49  8  7C  L;KM6  5:     input_general     Miscellaneous      �?      B�       A D� Q  A����        A����                         ��             0��    ��������             0��    ��������             0��    ��������             0��    ��������             0��    ��������             0��    �������� d   :�0�yE>10e-9��    �������� d   :�0�yE>10e-9��    ��������                            ����  ����:�0�yE>10e-9��d         ����  ����:�0�yE>10e-9��d   �     N  �����        d   :�0�yE>10e-9��    �������� d   :�0�yE>10e-9��    ��������1 Bit Inport1 Bit Inport                 ODigital<   Generic   ResetReset           ����  ��    �������� ����  ��    �������� ����  ��    �������� ����  ��    �������� ����  ��    �������� ����  ��    �������� ����  ��    ��������          ����            In F�    ����AA      INAA�>      Digital Instruments Generic                         `   `              `   �  �              `   �             �  `   `          �      11 �     I 11 �     O 11 �     � 11  D� O  R����       R����                          ��      x��    ��������      x��    ��������      x��    ��������      x��    ��������      x��    ��������      x��    �������� d   :�0�yE>10e-9��    �������� d   :�0�yE>10e-9��    ��������                            ����  ����:�0�yE>10e-9��d         ����  ����:�0�yE>10e-9��d   �     �   �����     ��   d   :�0�yE>10e-9��    �������� d   :�0�yE>10e-9��    ��������D� O  R����       R����                          ��      x��    ��������      x��    ��������      x��    ��������      x��    ��������      x��    ��������      x��    �������� d   :�0�yE>10e-9��    �������� d   :�0�yE>10e-9��    ��������                            ����  ����:�0�yE>10e-9��d         ����  ����:�0�yE>10e-9��d   �     �   �����     ��   d   :�0�yE>10e-9��    �������� d   :�0�yE>10e-9��    ��������OD� O  R����       R����                          ��      x��    ��������      x��    ��������      x��    ��������      x��    ��������      x��    ��������      x��    �������� d   :�0�yE>10e-9��    �������� d   :�0�yE>10e-9��    ��������                            ����  ����:�0�yE>10e-9��d         ����  ����:�0�yE>10e-9��d   �     ��       SJClkKRQQ' D� K  S����        S����                          ��      x��    ��������      x��    ��������      x��    ��������      x��    ��������      x��    ��������      x��    �������� d   :�0�yE>10e-9��    �������� d   :�0�yE>10e-9��    ��������                            ����  ����:�0�yE>10e-9��d         ����  ����:�0�yE>10e-9��d   �      W  �����     ��   d   :�0�yE>10e-9��    �������� d   :�0�yE>10e-9��    ��������D� L  J����       J����                          ��      x��    ��������      x��    ��������      x��    ��������      x��    ��������      x��    ��������      x��    �������� d   :�0�yE>10e-9��    �������� d   :�0�yE>10e-9��    ��������                             ����  ����:�0�yE>10e-9��d         ����  ����:�0�yE>10e-9��d   �     � W  �����     ��   d   :�0�yE>10e-9��    �������� d   :�0�yE>10e-9��    ��������D� M  Clk����       Clk����                          ��      x��    ��������      x��    ��������      x��    ��������      x��    ��������      x��    ��������      x��    �������� d   :�0�yE>10e-9��    �������� d   :�0�yE>10e-9��    ��������                            ����  ����:�0�yE>10e-9��d         ����  ����:�0�yE>10e-9��d   �     R W  �����     ��   d   :�0�yE>10e-9��    �������� d   :�0�yE>10e-9��    ��������D� N  K����       K����                          ��      x��    ��������      x��    ��������      x��    ��������      x��    ��������      x��    ��������      x��    �������� d   :�0�yE>10e-9��    �������� d   :�0�yE>10e-9��    ��������                            ����  ����:�0�yE>10e-9��d         ����  ����:�0�yE>10e-9��d   �     �	    �   \ 	 O 17 �   \ 	 � 17  D� Q  Q'����       Q'����                         �� �  :�0�ye>40ns��    ��������      x��    �������� �   I�����Z>25ns��    �������� �   I�����Z>25ns��    ��������      x��    �������� �   �?Y��K>13ns��    �������� d   :�0�yE>10e-9��    �������� d   :�0�yE>10e-9��    ��������                           ����  ����:�0�yE>10e-9��d         ����  ����:�0�yE>10e-9��d   �     \�   �����     ��  d   :�0�yE>10e-9��    �������� d   :�0�yE>10e-9��    ��������[	 17W  �����     ��   d   :�0�yE>10e-9��    �������� d   :�0�yE>10e-9��    ��������VD� P  Q����       Q����                         �� �  :�0�ye>40ns��    ��������      x��    �������� �   I�����Z>25ns��    �������� �   I�����Z>25ns��    ��������      x��    �������� �   �?Y��K>13ns��    �������� d   :�0�yE>10e-9��    �������� d   :�0�yE>10e-9��    ��������                            ����  ����:�0�yE>10e-9��d         ����  ����:�0�yE>10e-9��d   �     �    �   a  � 20 �    a   ��       _   @         _   @                 Output_Portc
�    �:   �  @   �-   �<   �  @   �,   h�5   �  �   i           g    f    �.   f�=   �  @   k                       �   port     �  �          Out4     !�                   ��                                                           @   port%�         �   `                   ����                                                 �   `   (�     @       @      ��                                                        #�    8       H                  ����
[negative]               ���                       8       H      8       H   >� (   ,   `   Q     ��                                                      (   ,   `   Q   (   ,   `   Q   [value]       �    �  �  (   ,   �   T   >�     $       <     ��                                                           $       <       $       <   [port.nbits]      <       ����            �      "Arial                    $       <   >�     ����j         ��                                                           ����j           ����j       	[refname]       �  h  �        �����       o  mpqrsn     Output_Port     Miscellaneous      �?      ��       port D� ����port����        port����                                         0��    ��������             0��    ��������             0��    ��������             0��    ��������             0��    ��������             0��    �������� d   :�0�yE>10e-9��    �������� d   :�0�yE>10e-9��    ��������                             ����  ����:�0�yE>10e-9��d         ����  ����:�0�yE>10e-9��d   �     at  �����     ��   d   :�0�yE>10e-9��    �������� d   :�0�yE>10e-9��    ��������Output_PortOutput_Port                 uDigital<   Generic   Out4Out4           ����  ��    �������� ����  ��    �������� ����  ��    �������� ����  ��    �������� ����  ��    �������� ����  ��    �������� ����  ��    ��������  ����    ����       ����  Out F�    ����portport       A �>      Digital Instruments Generic                                                                          lop                                 20  u` 20W  �����     ��   d   :�0�yE>10e-9��    �������� d   :�0�yE>10e-9��    ��������D� Q  Q'����       Q'����                         �� �  :�0�ye>40ns��    ��������      x��    �������� �   I�����Z>25ns��    �������� �   I�����Z>25ns��    ��������      x��    �������� �   �?Y��K>13ns��    �������� d   :�0�yE>10e-9��    �������� d   :�0�yE>10e-9��    ��������                           ����  ����:�0�yE>10e-9��d         ����  ����:�0�yE>10e-9��d   �     �    �   x  � 21  w 21W  �����     ��   d   :�0�yE>10e-9��    �������� d   :�0�yE>10e-9��    ��������109A/2 LS JK FF109A/2 LS JK FF / l             XYZ[V`wDigital<   Analog Devices   A5A5           ���� x��    �������� ���� x��    �������� �� hUMu�>30u��    �������� �r��b2U0*�C�-.6m��    �������� ���-C��6:�-.4m��    ��������  ������Mb�?8m��    ��������  Zb����Mbp?4m��    ��������          ����LS     2   :�0�y5>5n��    �������� ����    �xA33meg��    �������� �   I�����Z>25n��    �������� ,  ,i�)+`>30n��    ��������  �����     ��   d   :�0�yE>10e-9��    �������� d   :�0�yE>10e-9��    �������� 11�   �����     ��   d   :�0�yE>10e-9��    �������� d   :�0�yE>10e-9��    ��������D� P  Q����       Q����                         �� �  :�0�ye>40ns��    ��������      x��    �������� �   I�����Z>25ns��    �������� �   I�����Z>25ns��    ��������      x��    �������� �   �?Y��K>13ns��    �������� d   :�0�yE>10e-9��    �������� d   :�0�yE>10e-9��    ��������                            ����  ����:�0�yE>10e-9��d         ����  ����:�0�yE>10e-9��d   �     K �   �����        d   :�0�yE>10e-9��    �������� d   :�0�yE>10e-9��    ��������� 109A/2 LS JK FF109A/2 LS JK FF / l             � � � z� Digital<   Analog Devices   A1A1           ���� x��    �������� ���� x��    �������� �� hUMu�>30u��    �������� �r��b2U0*�C�-.6m��    �������� ���-C��6:�-.4m��    ��������  ������Mb�?8m��    ��������  Zb����Mbp?4m��    ��������    `     ����LS     2   :�0�y5>5n��    �������� ����    �xA33meg��    �������� �   I�����Z>25n��    �������� ,  ,i�)+`>30n��    ��������  �����         d   :�0�yE>10e-9��    �������� d   :�0�yE>10e-9��    ���������  13�   �����     ��   d   :�0�yE>10e-9��    �������� d   :�0�yE>10e-9��    ��������TD� P  Q����       Q����                         �� �  :�0�ye>40ns��    ��������      x��    �������� �   I�����Z>25ns��    �������� �   I�����Z>25ns��    ��������      x��    �������� �   �?Y��K>13ns��    �������� d   :�0�yE>10e-9��    �������� d   :�0�yE>10e-9��    ��������                            ����  ����:�0�yE>10e-9��d         ����  ����:�0�yE>10e-9��d   �     K �   �����     ��  d   :�0�yE>10e-9��    �������� d   :�0�yE>10e-9��    ��������� 109A/2 LS JK FF109A/2 LS JK FF / l             � � � � T{� Digital<   Analog Devices   A2A2           ���� x��    �������� ���� x��    �������� �� hUMu�>30u��    �������� �r��b2U0*�C�-.6m��    �������� ���-C��6:�-.4m��    ��������  ������Mb�?8m��    ��������  Zb����Mbp?4m��    ��������          ����LS     2   :�0�y5>5n��    �������� ����    �xA33meg��    �������� �   I�����Z>25n��    �������� ,  ,i�)+`>30n��    ��������  �����     ��  d   :�0�yE>10e-9��    �������� d   :�0�yE>10e-9��    ���������  7�   �����     ��   d   :�0�yE>10e-9��    �������� d   :�0�yE>10e-9��    ��������U� _109A/2 LS JK FF109A/2 LS JK FF / l             � � � � U� _Digital<   Analog Devices   A3A3           ���� x��    �������� ���� x��    �������� �� hUMu�>30u��    �������� �r��b2U0*�C�-.6m��    �������� ���-C��6:�-.4m��    ��������  ������Mb�?8m��    ��������  Zb����Mbp?4m��    ��������          ����LS     2   :�0�y5>5n��    �������� ����    �xA33meg��    �������� �   I�����Z>25n��    �������� ,  ,i�)+`>30n��    ��������  �����     ��  d   :�0�yE>10e-9��    �������� d   :�0�yE>10e-9��    ��������Y 16  � 16 � ^Sby
�              S   
�   �       �  J   
�   l       @  Clk    
�   �3   `  �   �1   �   �  �   � 	      �     	            �  K    
�   3     `  R   
�   j  @  �  Q   
�   �6   �  �             @  �  Q'    `  �          A5     !�                    ��                                                       `   `   S!�                   ��                                                          �   J!�                   ��                                                          �   Clk!�                   ��                                                          �   K!�                   ��                                                      `      R!�                   ��                                                      �   �   Q!�                   ��                                                      �   �   Q'%�     �   �                     ����                                             �   �      (� `   `   `   p     ��                                                        (�     �       �    	 ��        	                                                (�     �       �    
 ��        
                                                (�     �      �     ��                                                        (� �   �   �   �     ��                                                        (� �   �   �   �     ��                                                        (� (   �       �     ��                                                        (�     �   (   �     ��                                                        (� `     `        ��                                                        #� X   p   h   �                  �                                           X   p   h   �   X   p   h   �   #� X      h                    �                                           X      h     X      h     #�    �       �                  �                                              �       �      �       �   #� �   �   �   �                  �                                           �   �   �   �   �   �   �   �   >� (   �   0   �     ��                                                      (   �   0   �   (   �   0   �   j       �  �  �  &  (   �   \   �   >� 4   �   \   �     ��                                                      4   �   \   �   4   �   \   �   clk       �  �  t  �  4   �   h   �   >� (   �   8   �     ��                                                      (   �   8   �   (   �   8   �   k       �  P    �  (   �   \   �   >�     0   b   X     ��                                                           0   b   X       0   b   X   	[refname]       �  p  �        0   �   T   >�        �   0     ��                                                              �   0          �   0   	[devname]        ����������������       �   0   ! �����������������      �  �������      �     74109/2    74109/2 IEEEMiscellaneous      �?    /  W  A F�    ����SS      INAS ���    F�   ����JJ      INAJE>1   F�   ����ClkClk      INAClk>10   F�   ����KK      INAK       F�   ����RR      INAR>�    F�   ����QQ      OUTAQ���    F�   ����Q'Q'      TRIAQ'� d   F�    ����SS      INBS�       F�   ����JJ      INBJ�     F�   ����ClkClk      INBClk       F�   ����KK      INBKA�>    F�   ����RR      INBR����   F�   ����QQ      OUTBQ�     F�   ����Q'Q'      TRIBQ'�     
Flip Flops2JK pos edge triggered flip-flop w/preset and clearGenericDO16             3  � � � Z 3  O 3 � R� ]
�              S    
�   �   �  �   �    �-   `  �   �&   �.   `  @   �   	     �    �%   �   @  �   �   �      �   ��#   ��+   �
  �   ��   �   �	  �   �        �    �$   �,   �
  @   �        �                   �    �       �    �    �    �   ��*   �  �   �                     �  J    
�   f       @  Clk    
�   �   �  �   �   �    @  �   �       �                 �  K    
�   /     `  R    
�   �   @  �  Q    
�   �  @  �  Q'     �  �          A3     !�                    ��                                                       `   `   S!�                   ��                                                          �   J!�                   ��                                                          �   Clk!�                   ��                                                          �   K!�                   ��                                                      `      R!�                   ��                                                      �   �   Q!�                   ��                                                      �   �   Q'%�     �   �                     ����                                             �   �      (� `   `   `   p     ��                                                        (�     �       �    	 ��        	                                                (�     �       �    
 ��        
                                                (�     �      �     ��                                                        (� �   �   �   �     ��                                                        (� �   �   �   �     ��                                                        (� (   �       �     ��                                                        (�     �   (   �     ��                                                        (� `     `        ��                                                        #� X   p   h   �                  �                                           X   p   h   �   X   p   h   �   #� X      h                    �                                           X      h     X      h     #�    �       �                  �                                              �       �      �       �   #� �   �   �   �                  �                                           �   �   �   �   �   �   �   �   >� (   �   0   �     ��                                                      (   �   0   �   (   �   0   �   j       �  �    &  (   �   \   �   >� 4   �   \   �     ��                                                      4   �   \   �   4   �   \   �   clk         �  �  �  4   �   h   �   >� (   �   8   �     ��                                                      (   �   8   �   (   �   8   �   k       �  P  (  �  (   �   \   �   >�     0   b   X     ��                                                           0   b   X       0   b   X   	[refname]       �  p  �        0   �   T   >�        �   0     ��                                                              �   0          �   0   	[devname]        ����������������       �   0   ! �����������������      �  �������      �     74109/2    74109/2 IEEEMiscellaneous      �?    /  �   A F�    ����SS      INAS�0�    F�   ����JJ      INAJyE>   F�   ����ClkClk      INAClk   �   F�   ����KK      INAK       F�   ����RR      INAR      F�   ����QQ      OUTAQzzzz   F�   ����Q'Q'      TRIAQ'�     F�    ����SS      INBS        F�   ����JJ      INBJ 0�   F�   ����ClkClk      INBClk      F�   ����KK      INBK�
    F�   ����RR      INBR      F�   ����QQ      OUTBQ       F�   ����Q'Q'      TRIBQ'����   
Flip Flops2JK pos edge triggered flip-flop w/preset and clearGenericDO16              12 �    K    ��       _   @         _   @                 Output_Port�
�    �       �   port     �
  �          Out1     !�                   ��                                                           @   port%�         �   `                   ����                                                 �   `   (�     @       @      ��    ����                                                #�    8       H                  ����
[negative]               ���                       8       H      8       H   >� (   ,   E   Q     ��                                                      (   ,   E   Q   (   ,   E   Q   [value]       �
    P  �  (   ,   �   T   >�     $       <     ��                                                           $       <       $       <   [port.nbits]      <       ����            �      "Arial                    $       <   >�     ����j         ��                                                           ����j           ����j       	[refname]       �
  h  �        �����       �  ������     Output_Port     Miscellaneous      �?      ��       port D� ����port����        port����                                         0��    ��������             0��    ��������             0��    ��������             0��    ��������             0��    ��������             0��    �������� d   :�0�yE>10e-9��    �������� d   :�0�yE>10e-9��    ��������                             ����  ����:�0�yE>10e-9��d         ����  ����:�0�yE>10e-9��d   �     K �  �����     ��   d   :�0�yE>10e-9��    �������� d   :�0�yE>10e-9��    ��������Output_PortOutput_Port                 �Digital<   Generic   Out1Out1           ����  ��    �������� ����  ��    �������� ����  ��    �������� ����  ��    �������� ����  ��    �������� ����  ��    �������� ����  ��    ��������          ����       ����  Out F�    ����portport       A �>      Digital Instruments Generic                                                                                                              12 �    K    ��	       _   @         _   @                 Output_Port�
�    �       �   port     `  �          Out2     !�                   ��                                                           @   port%�         �   `                   ����                                                 �   `   (�     @       @      ��    ����                                                #�    8       H                  ����
[negative]               ���                       8       H      8       H   >� (   ,   E   Q     ��                                                      (   ,   E   Q   (   ,   E   Q   [value]       �    0  �  (   ,   �   T   >�     $       <     ��                                                           $       <       $       <   [port.nbits]      <       ����            �      "Arial                    $       <   >�     ����j         ��                                                           ����j           ����j       	[refname]       �  h  �        �����              Output_Port     Miscellaneous      �?      ��       port D� ����port����        port����                                         0��    ��������             0��    ��������             0��    ��������             0��    ��������             0��    ��������             0��    �������� d   :�0�yE>10e-9��    �������� d   :�0�yE>10e-9��    ��������                             ����  ����:�0�yE>10e-9��d         ����  ����:�0�yE>10e-9��d   �     K 	  �����     ��   d   :�0�yE>10e-9��    �������� d   :�0�yE>10e-9��    ��������Output_PortOutput_Port                 
Digital<   Generic   Out2Out2           ����  ��    �������� ����  ��    �������� ����  ��    �������� ����  ��    �������� ����  ��    �������� ����  ��    �������� ����  ��    ��������         ����       ����  Out F�    ����portport       A �>      Digital Instruments Generic                                                                                                              12  �
z� {�  12  I 12 � � QM � 
�              S    
�   �      �  J   
�   `       @  Clk   
�   �      �   �"   �   �	  �                            �  K   
�   +     `  R   
�   �  @  �  Q   
�   �  @  �  Q'       �          A2     !�                    ��                                                       `   `   S!�                   ��                                                          �   J!�                   ��                                                          �   Clk!�                   ��                                                          �   K!�                   ��                                                      `      R!�                   ��                                                      �   �   Q!�                   ��                                                      �   �   Q'%�     �   �                     ����                                             �   �      (� `   `   `   p     ��    ? �                                                (�     �       �    	 ��        	                                                (�     �       �    
 ��    � �
                                                (�     �      �     ��    ����                                                (� �   �   �   �     ��                                                        (� �   �   �   �     ��                                                        (� (   �       �     ��                                                        (�     �   (   �     ��                                                        (� `     `        ��                                                        #� X   p   h   �                  �                                           X   p   h   �   X   p   h   �   #� X      h                    �                                           X      h     X      h     #�    �       �                  �                                              �       �      �       �   #� �   �   �   �                  �                                           �   �   �   �   �   �   �   �   >� (   �   0   �     ��                                                      (   �   0   �   (   �   0   �   j       x  �  �  &  (   �   \   �   >� 4   �   \   �     ��                                                      4   �   \   �   4   �   \   �   clk       �  �    �  4   �   h   �   >� (   �   8   �     ��                                                      (   �   8   �   (   �   8   �   k       x  P  �  �  (   �   \   �   >�     0   b   X     ��                                                           0   b   X       0   b   X   	[refname]       `  p  (        0   �   T   >�        �   0     ��                                                              �   0          �   0   	[devname]        ����������������       �   0   !  !"#+,-      %  '(./)*$      &     74109/2    74109/2 IEEEMiscellaneous      �?    /  �   A F�    ����SS      INAS @    F�   ����JJ      INAJ ��   F�   ����ClkClk      INAClk��u�   F�   ����KK      INAK����   F�   ����RR      INAR  ��   F�   ����QQ      OUTAQ      F�   ����Q'Q'      TRIAQ'� x   F�    ����SS      INBS        F�   ����JJ      INBJ����   F�   ����ClkClk      INBClk  ��   F�   ����KK      INBKx'    F�   ����RR      INBRtrue   F�   ����QQ      OUTBQ ��   F�   ����Q'Q'      TRIBQ'��u�   
Flip Flops2JK pos edge triggered flip-flop w/preset and clearGenericDO16             14 P �  � � � E X  14  �� 14 � S � L � 
�              S    
�   �       �  J   
�   r       @  Clk   
�         �  K   
�   '     `  R   
�   �  @  �  Q   
�     @  �  Q'    �  �          A1     !�                    ��                                                       `   `   S!�                   ��                                                          �   J!�                   ��                                                          �   Clk!�                   ��                                                          �   K!�                   ��                                                      `      R!�                   ��                                                      �   �   Q!�                   ��                                                      �   �   Q'%�     �   �                     ����                                             �   �      (� `   `   `   p     ��    t �                                                (�     �       �    	 ��    ����	                                                (�     �       �    
 ��       
                                                (�     �      �     ��    ����                                                (� �   �   �   �     ��    ����                                                (� �   �   �   �     ��    ����                                                (� (   �       �     ��    ����                                                (�     �   (   �     ��    -9 �                                                (� `     `        ��                                                       #� X   p   h   �                  �                                           X   p   h   �   X   p   h   �   #� X      h                    �                                           X      h     X      h     #�    �       �                  �                                              �       �      �       �   #� �   �   �   �                  �                                           �   �   �   �   �   �   �   �   >� (   �   0   �     ��                                                      (   �   0   �   (   �   0   �   j       �  �    &  (   �   \   �   >� 4   �   \   �     ��                                                      4   �   \   �   4   �   \   �   clk         �  �  �  4   �   h   �   >� (   �   8   �     ��                                                      (   �   8   �   (   �   8   �   k       �  P  (  �  (   �   \   �   >�     0   b   X     ��                                                           0   b   X       0   b   X   	[refname]       �  p  �        0   �   T   >�        �   0     ��                                                              �   0          �   0   	[devname]        ����������������       �   0   ! EFGHIJKLMNOPQRZ[\      T  VW]^XYS      U4     74109/2    74109/2 IEEEMiscellaneous      �?    /  �   A F�    ����SS      INASield    F�   ����JJ      INAJ       F�   ����ClkClk      INAClk      F�   ����KK      INAK  �   F�   ����RR      INAR      F�   ����QQ      OUTAQ      F�   ����Q'Q'      TRIAQ'���:   F�    ����SS      INBS�0�    F�   ����JJ      INBJx��    F�   ����ClkClk      INBClk       F�   ����KK      INBK       F�   ����RR      INBR  �    F�   ����QQ      OUTBQ�    F�   ����Q'Q'      TRIBQ' �     
Flip Flops2JK pos edge triggered flip-flop w/preset and clearGenericDO16              I O � V � 	 !� � � d    � R � K � � � \� � � ax5 5 5 0m � k i _ g c ] a [ � Y o � q � .   $&(  *���e ��,���� � � 2igk� � �   A A A ��'� �   �` l +��  �f �/� �� ^ � p r X d \ b Z     # %)-������ � � �3j�h j n f1hl�                 
 ��@ ����        ����������             0     ���������� ����      @5     ����������  ʚ;�������?.1     ����������@ ����       ���������� ����       ���������� ����       ���������� ����       ���������� ���� true
     ���������� ����  false     ��������               
                  �� ����        ���������� ����       ����������  ����       ����������@ ����       ����������@ ����       ��������               
                  �� ����        ���������� ����       ����������@ ����       ����������  ����       ���������� ����       ���������� ����       ���������� ����       ���������� ����       ���������� ����       ���������� ����       ���������� ����       ��������               
                 �� ����dec     ���������� ����     @�@1k     ���������� ����    ��.A1meg     ���������� ����       20     ���������� ���� true     ���������� ���� true     ���������� ���� true	     ���������� ����  false
     ��������               
                 ��  ����        ����������  ����       ����������  ����       ���������� ����dec     ���������� ����       ���������� ����       ���������� ����  	     ���������� ����  
     ��������               
                  	 �� ����        ���������� ����       ���������� ����       ���������� ����       ���������� ����       ���������� ����       ���������� ����       ���������� ����       ���������� ����       ��������               
                 �� ����        ���������� ����       ���������� ����       ���������� ����dec     ���������� ����       ��������               
                     ��             0      ���������� ��� ����MbP?1m     ���������� �� �h㈵��>10u     ���������� '  ���ư>1u     ���������� ���� true     ���������� ����  false     ���������� ���� true     ���������� ����  false     ��������               
                 �� ����     @�@1K      ����������  ����       ����������  ����       ����������  ����       ��������               
         ��              ��  ����        ��������              
                  ��  ����        ��������              
                                  
                 ��@ ����        ����������@ ����       ���������� ����       ���������� ����       ���������� ����       ���������� ����       ���������� ����       ���������� ����       ���������� ����       ���������� ���� true	     ���������� ����  false
     ���������� ���� true     ���������� ����  false     ��������               
                 �� ����       5      ���������� ����       5     ���������� ����       5     ���������� ����       5     ���������� ����       ���������� ����  	     ���������� ����  
     ���������� ����       ���������� ����       ���������� ����       ���������� ���� true     ����������@ ����       ����������@ ����       ���������� ����       ���������� ����       ���������� ����       ���������� ����dec     ���������� ����       ���������� ����       ���������� ����       ���������� ���� true     ���������� ���� true     ���������� ���� true     ���������� ����  false     ���������� ���� true     ���������� ����  false      ���������� ���� true!     ���������� ����  false"     ��������               
                        �� ����       5      ���������� ����       5     ���������� ����       5     ���������� ����       5     ���������� ����       ���������� ����  	     ���������� ����  
     ���������� ����       ���������� ����       ���������� ����       ���������� ���� true     ����������@ ����       ����������@ ����       ���������� ����       ���������� ����       ���������� ����       ���������� ����dec     ���������� ����       ���������� ����       ���������� ����       ���������� ���� true     ���������� ���� true     ���������� ���� true     ���������� ����  false     ���������� ���� true     ���������� ����  false      ���������� ���� true!     ���������� ����  false"     ��������               
                 �� ����       5      ���������� ����       5     ���������� ����       5     ���������� ����       5     ���������� ����       ���������� ����  	     ���������� ����  
     ���������� ����       ���������� ����       ���������� ����       ���������� ���� true     ����������@ ����       ����������@ ����       ���������� ����       ���������� ����       ���������� ����       ���������� ����dec     ���������� ����       ���������� ����       ���������� ����       ���������� ���� true     ���������� ���� true     ���������� ���� true     ���������� ����  false     ���������� ���� true     ���������� ����  false      ���������� ���� true!     ���������� ����  false"     ��������               
                 �� ����       5      ���������� ����       5     ���������� ����       5     ���������� ����       5     ���������� ����       ���������� ����  	     ���������� ����  
     ���������� ����       ���������� ����       ���������� ����       ���������� ���� true     ����������@ ����       ����������@ ����       ���������� ����       ���������� ����       ���������� ����       ���������� ����dec     ���������� ����       ���������� ����       ���������� ����       ���������� ���� true     ���������� ���� true     ���������� ���� true     ���������� ����  false     ���������� ���� true     ���������� ����  false      ���������� ���� true!     ���������� ����  false"     ��������               
                 ��@ ����        ����������@ ����       ���������� ����       ���������� ����       ���������� ����       ���������� ����       ���������� ����       ���������� ����       ���������� ����decade     ���������� ���� true     ���������� ���� true     ���������� ���� true     ���������� ����  false     ��������               
                 �� ����        ���������� ����       ����������@ ����       ����������  ����       ���������� ����       ���������� ����       ���������� ����       ���������� ����       ���������� ����       ���������� ����       ���������� ����       ��������               
                        �� ����dec     ���������� ����     @�@1k     ���������� ����    ��.A1meg     ���������� ����       20     ���������� ����        0     ���������� ����        0     ���������� ���� true	     ���������� ���� true
     ���������� ����      I@50     ���������� ���� true     ���������� ����  false     ��������               
                          / �� ���� x'     ����������     �-���q=1E-12     ���������� @B -C��6?1E-4     ���������� ���� x     ���������� ���� x     ���������� ���� x     ���������� ���� x     ���������� ���� x     ���������� ���� x     ���������� ���� x	     ���������� ���� x!     ���������� ����    �  500
     ���������� ���� x     ���������� ����    �  500     ���������� ���� x$     ���������� ���� x$     ���������� ���� x%     ���������� ���� x"     ����������  ���� x*     ���������� ���� x     ���������� ���� x     ���������� ���� x     ���������� ���� x&     ���������� ���� x     ���������� ���� x     ���������� ���� x     ���������� ���� x+     ���������� ���� x,     ���������� ���� x-     ���������� ���� xg     ���������� ���� xf     ���������� ���� xd     ���������� ���� xe     ���������� ���� xh     ���������� ���� xj     ���������� ���� xi     ���������� ���� xk     ���������� ����    e��A1Gl     ����������             0�     ���������� ����      @5�     ���������� ����      @2.5�     ���������� ����      �?.5�     ���������� ����      @4.5�     ���������� 
   ��&�.>1n�     ���������� 
   ��&�.>1n�     ���������� 
   ��&�.>1n�     ���������� 
   ��&�.>1n�     ��������                                  Ariald        ��=i|�x�  �=i,� ��/i    ��=i|�x�  �=i,� ��/i ��  COpAnal                         
                        ����                                   ��=i|�x�  �=i,� ��/i    ��=i|�x�  �=i,� ��/i ��  CDCsweep       
 mnopqrstuv               
                      ����                                   ��=i|�x�  �=i,� ��/i    ��=i|�x�  �=i,� ��/i ��  CACsweep        ��������               
                      ����                                  ��=i|�x�  �=i,� ��/i    ��=i|�x�  �=i,� ��/i �� 
 CTranSweep        ��������               
                      ����                                   ��=i|�x�  �=i,� ��/i    ��=i|�x�  �=i,� ��/i ��  CACdisto        �����               
                          ����                                  ��=i|�x�  �=i,� ��/i    ��=i|�x�  �=i,� ��/i ��        �� ����        ���������� ����       ���������� ����       ���������� ����dec     ���������� ����       ��������               
         �                ����                                  ��=i|�x�  �=i,� ��/i    ��=i|�x�  �=i,� ��/i ��        �� ����        ���������� ����       ���������� ����       ���������� ����dec     ���������� ����       ��������               
         �                ����                                  ��=i|�x�  �=i,� ��/i    ��=i|�x�  �=i,� ��/i ��        �� ����        ���������� ����       ���������� ����       ���������� ����dec     ���������� ����       ��������               
         d                ����                                  ��=i|�x�  �=i,� ��/i    ��=i|�x�  �=i,� ��/i ��        �� ����        ���������� ����       ���������� ����       ���������� ����dec     ���������� ����       ��������               
                          ����                                  ��=i|�x�  �=i,� ��/i    ��=i|�x�  �=i,� ��/i ��        �� ����        ���������� ����       ���������� ����       ���������� ����dec     ���������� ����       ��������               
         �            	    ����                                  ��=i|�x�  �=i,� ��/i    ��=i|�x�  �=i,� ��/i ��  CACnoise        ��������               
                   
    ����            �                   ��=i|�x�  �=i,� ��/i    ��=i|�x�  �=i,� ��/i ��                        
                        ����           ����                   ��=i|�x�  �=i,� ��/i    ��=i|�x�  �=i,� ��/i ��  CFourier        ����               
         ��                  ����            ����                   ��=i|�x�  �=i,� ��/i    ��=i|�x�  �=i,� ��/i ��  CACpz        	 ���������               
                       ����                                   ��=i|�x�  �=i,� ��/i    ��=i|�x�  �=i,� ��/i ��  CDCtf         wxyz{               
                       ����                                  ��=i|�x�  �=i,� ��/i    ��=i|�x�  �=i,� ��/i ��  CDCsens         |}~�������               
                       ����            �� �                   ��=i|�x�  �=i,� ��/i    ��=i|�x�  �=i,� ��/i                 ����            ����                   ��=i|�x�  �=i,� ��/i    ��=i|�x�  �=i,� ��/i ��  CShow         �              
                       ����            ����                   ��=i|�x�  �=i,� ��/i    ��=i|�x�  �=i,� ��/i ��  CShowmod         �              
                       ����                                   ��=i|�x�  �=i,� ��/i    ��=i|�x�  �=i,� ��/i �� 
 CLinearize        ��  ����        ��������               
                      ����                                  ��=i|�x�  �=i,� ��/i    ��=i|�x�  �=i,� ��/i ��  CParamTranSweep        �������������               
                      ����            ls �                   ��=i|�x�  �=i,� ��/i    ��=i|�x�  �=i,� ��/i �             ����            #� �                   ��=i|�x�  �=i,� ��/i    ��=i|�x�  �=i,� ��/i ��  CParamACSweep        0123456789:;<               
                      ����           ����                   ��=i|�x�  �=i,� ��/i    ��=i|�x�  �=i,� ��/i ��  CMonteCarlo_op        ����������������������������               
                             ����            ����                   ��=i|�x�  �=i,� ��/i    ��=i|�x�  �=i,� ��/i ��  CMonteCarlo_dc        ����������������������������               
                      ����                                   ��=i|�x�  �=i,� ��/i    ��=i|�x�  �=i,� ��/i ��  CMonteCarlo_ac        �������� 	
               
                      ����                                 ��=i|�x�  �=i,� ��/i    ��=i|�x�  �=i,� ��/i ��  CMonteCarlo_tran         !"#$%&'()*+,-./               
                      ����            �  �                   ��=i|�x�  �=i,� ��/i    ��=i|�x�  �=i,� ��/i ��  CACsens        =>?@ABCDEFG               
                             ����           ����                   ��=i|�x�  �=i,� ��/i    ��=i|�x�  �=i,� ��/i ��  CNetworkAnalysis        HIJKLMNOPQR               
                      ����           ����                   ��=i|�x�  �=i,� ��/i    ��=i|�x�  �=i,� ��/i                 ����                                 >           ��   CDigSimResTemplate    	   ��   TDigitalSignal            Set       ����                        ΃            U1        ����                        ΃            In2        ����                        ΃            Out1        ����                        ΃            Out2        ����                        ΃            Out3        ����                        ΃            Reset        ����                        ΃            Out4        ����                                  ���       ����  ����:�0�yU>+20.00n���   ����                       Arial����                       Arial����                       Arial                                          ����  ����        0��          ����  ����        0��                     �               ����  �����       200������          0.000000e+000��    ��������      0.000000e+000��    ��������      0.000000e+000��    ��������   ����                       Arial����                       Arial����                       Arial����                       Arial                        �     �   �  �                     ����  ��    ��������   A  DO16�16 pin small outline package                                                                                                                                                                                                                              ����   ��   CPackageAliasSuperPCBStandardSO16      ׃EagleBURR.LBRSO16-1      ׃Orcad SOG.050/16/WG.255/L.400      ׃Pads SO16NB      ׃	UltiboardL7IC.l55$SO16      ׃Eaglesmd-ipc.lbrSO16             A                A  DO16�16 pin small outline package                                                                                                                                                                                                                              ����   ������        B                A  DO16�16 pin small outline package                                                                                                                                                                                                                              ����   ������        A                                              @  DO14�14 pin small outline package                                                                                                                                                                                                                              ����   ׃SuperPCBStandardSO14      ׃EagleBURR.LBRSO14      ׃Orcad SOG.050/14/WG.244/L.350      ׃Pads SO14NB      ׃	UltiboardL7IC.l55$SO14      ׃Eagleburr-brown.lbrSO14             A                                                                  A  DO16�16 pin small outline package                                                                                                                                                                                                                              ����   ������        B                          �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                   ط�     ����t� ؙ�     <�     N   N   ��     ؙ� N                  2         �                 � � �           k t     ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                   ط�     ����t� ؙ�     <�     N   N   ��     ؙ� N                  2         �                 � � �           k t     ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                   ط�     ����t� ؙ�     <�     N   N   ��     ؙ� N                  2         �                 � � �           k t     ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                   ط�     ����t� ؙ�     <�     N   N   ��     ؙ� N                  2         �                 � � �           k t     ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                   ط�     ����t� ؙ�     <�     N   N   ��     ؙ� N                  2         �                 � � �           k t     ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                   ط�     ����t� ؙ�     <�     N   N   ��     ؙ� N                  2         �                 � � �           k t     ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                   ط�     ����t� ؙ�     <�     N   N   ��     ؙ� N                  2         �                 � � �           k t     ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                   ط�     ����t� ؙ�     <�     N   N   ��     ؙ� N                  2         �                 � � �           k t     ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                   ط�     ����t� ؙ�     <�     N   N   ��     ؙ� N                  2         �                 � � �           k t     ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                   ط�     ����t� ؙ�     <�     N   N   ��     ؙ� N                  2         �                 � � �           k t     ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                   ط�     ����t� ؙ�     <�     N   N   ��     ؙ� N                  2         �                 � � �           k t     ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                   ط�     ����t� ؙ�     <�     N   N   ��     ؙ� N                  2         �                 � � �           k t     ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                   ط�     ����t� ؙ�     <�     N   N   ��     ؙ� N                  2         �                 � � �           k t     ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                   ط�     ����t� ؙ�     <�     N   N   ��     ؙ� N                  2         �                 � � �           k t     ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                   ط�     ����t� ؙ�     <�     N   N   ��     ؙ� N                  2         �                 � � �           k t     ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                   ط�     ����t� ؙ�     <�     N   N   ��     ؙ� N                  2         �                 � � �           k t     ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                   ط�     ����t� ؙ�     <�     N   N   ��     ؙ� N                  2         �                 � � �           k t     ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                   ط�     ����t� ؙ�     <�     N   N   ��     ؙ� N                  2         �                 � � �           k t     ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                   ط�     ����t� ؙ�     <�     N   N   ��     ؙ� N                  2         �                 � � �           k t     ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                   ط�     ����t� ؙ�     <�     N   N   ��     ؙ� N                  2         �                 � � �           k t     ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                   ط�     ����t� ؙ�     <�     N   N   ��     ؙ� N                  2         �                 � � �           k t     ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                   ط�     ����t� ؙ�     <�     N   N   ��     ؙ� N                  2         �                 � � �           k t     ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                   ط�     ����t� ؙ�     <�     N   N   ��     ؙ� N                  2         �                 � � �           k t     ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                   ط�     ����t� ؙ�     <�     N   N   ��     ؙ� N                  2         �                 � � �           k t     ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                   ط�     ����t� ؙ�     <�     N   N   ��     ؙ� N                  2         �                 � � �           k t     ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                   ط�     ����t� ؙ�     <�     N   N   ��     ؙ� N                  2         �                 � � �           k t     ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                   ط�     ����t� ؙ�     <�     N   N   ��     ؙ� N                  2         �                 � � �           k t     ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                   ط�     ����t� ؙ�     <�     N   N   ��     ؙ� N                  2         �                 � � �           k t     ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                   ط�     ����t� ؙ�     <�     N   N   ��     ؙ� N                  2         �                 � � �           k t     ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                   ط�     ����t� ؙ�     <�     N   N   ��     ؙ� N                  2         �                 � � �           k t     ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                               �� 	 CTitleBox                        ��=i    ����                  �	                  %�         �  @                  ���                                                  �  @  (�     <   �  <     ��    D��                                                (�     |   �  |     ��       �                                                (�     �   �  �     ��    ��                                                (�     �   �  �     ��    �@�                                                >� h      t  4     ��                                                      h      t  4   h      t  4   [title]                                       >� �   H   �  x     ��                                                      �   H   �  x   �   H   �  x   [description]                                       >� P   �   X  �     ��                                                      P   �   X  �   P   �   X  �   [id]                                       >� �   �   �  �     ��                                                      �   �   �  �   �   �   �  �   
[designer]                                       >�      ]   1    ��        	                                                   ]   1       ]   1  Date :       �  4  �  �                  >� p     x  4   	 ��        
                                              p     x  4  p     x  4  [date]                                       >�       U   1    
 ��                                                            U   1         U   1   Title :       �  4  �  �                  >�    L   �   q     ��                                                         L   �   q      L   �   q   Description :       �  �  �   �                  >�    �   8   �     ��                                                         �   8   �      �   8   �   ID :       �  �  8  J                  >�    �   �   �     ��                                                         �   �   �      �   �   �   
Designer :       �  t  p   
                   ��������������          �     	title box     Miscellaneous      �?    9 
 ��  CParamSubBehavior    
 ��  ����        ����������  ����       ����������  ����       ����������  ����       ����������  ����       ����������  ����       ����������  ����       ����������  ����       ����������  ����       ����������  ����  	     ��������        9                      �               ������   CParamSubModelType�� ����  
   ��  	 CParmDefn            title                �            description                �            id                �            designer                �            Date :                �            date                �            Title :                �            Description :                �            ID :                �            
Designer :                            ����             `         �?�� 	 CGraphDoc�  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                   ��t�u��t�	u����t �t �tp�t,�t�t�u u8�t�u             2         �                 � � �           @�t    ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                         �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                   ��t�u��t�	u����t �t        ,�t�t�u          u        ΃            In1        ����                        ΃            U1        ����                        ΃            In2        ����                        ΃            In3        ����                        ΃            Out1        ����                        ΃            Out2        ����                        ΃            Out3        ����                            2         �                 � � �                   ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                        ��SetU1In2Out1Out2Out3ResetOut4                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                     1m  0                            100   100                                                           1m  0                            100   100                              1m  0                            100   100                              1m  0                            100   100                                                 
               1m  0                            100   100                            ��   CPartPackage�t� ��   CPackageA  DO16�16 pin small outline package                                                                                                                                                                                                                              ����   ������   ��t�    ���� �@  DO14�14 pin small outline package                                                                                                                                                                                                                              ����   ������    ��   CMiniPartPin    ����SS     INS�      �   ����JJ     INJ�     �   ����ClkClk     INClk�     �   ����KK     INK�     �   ����RR     INR�     �   ����QQ     OUTQ�     �   ����Q'Q'     TRIQ'�       I   ��   CPackagePin 2 J   A1J&� 3 K   A~1K&� 4 Clk   A1CLK&� 5 S   A~1PR&� 1 R   A~1CLR&� 6 Q   A1Q&� 7 Q'   A~1Q&� 8  GND  COMGND&� 9 Q'  	 B~2Q&� 10 Q  
 B2Q&� 11 S   B~2PR&� 12 Clk   B2CLK&� 13 K   B~2K&� 14 J   B2J&� 15 R   B~2CLR&� 16  VCC  COMVCC2JK pos edge triggered flip-flop w/preset and clear
Flip FlopsGenericC      74109 A74LS109DA1               DIP1674LS109D74LS109D��  CXSpiceBehavior       jkclksetresetoutNout ��   CBehPin I  j����    �  j����                         ��9� I  k����   �  k����                         ��9� I  clk����   �  clk����                         ��9� I  set����   �  set����                         ��9� I  reset����   �  reset����                         ��9� I  out����   �  out����                        ��9� I  Nout����   �  Nout����                        ��74LS109A (Xspice)74LS109A (Xspice)  8               :;<=>?@Digital<   Generic                       * time value jJkKresetRoutQsetSclkClkNoutQ' JjKkQ'NoutQoutRresetClkclkSset                                                              �    ����SS     INS�      �   ����JJ     INJ�     �   ����ClkClk     INClk�     �   ����KK     INK�     �   ����RR     INR�     �   ����QQ     OUTQ�     �   ����Q'Q'     TRIQ'�       I   '()*+,-./01234562JK pos edge triggered flip-flop w/preset and clear
Flip FlopsGenericC      74109 A74LS109DA1               DIP1674LS109D74LS109D7�       jkclksetresetoutNout 9� I  j����    �  j����                         ��9� I  k����   �  k����                         ��9� I  clk����   �  clk����                         ��9� I  set����   �  set����                         ��9� I  reset����   �  reset����                         ��9� I  out����   �  out����                        ��9� I  Nout����   �  Nout����                        ��74LS109A (Xspice)74LS109A (Xspice)  8               IJKLMNODigital<   Generic                       * time value jJkKresetRoutQsetSclkClkNoutQ' JjKkQ'NoutQoutRresetClkclkSset                                                              �    ����SS     INS�      �   ����JJ     INJ�     �   ����ClkClk     INClk�     �   ����KK     INK�     �   ����RR     INR�     �   ����QQ     OUTQ�     �   ����Q'Q'     TRIQ'�      O �   &� 2 J   A1J&� 3 K   A~1K&� 4 Clk   A1CLK&� 5 S   A~1PR&� 1 R   A~1CLR&� 6 Q   A1Q&� 7 Q'   A~1Q&� 8  GND  COMGND&� 9 Q'  	 B~2Q&� 10 Q  
 B2Q&� 11 S   B~2PR&� 12 Clk   B2CLK&� 13 K   B~2K&� 14 J   B2J&� 15 R   B~2CLR&� 16  VCC  COMVCC2JK pos edge triggered flip-flop w/preset and clear
Flip FlopsGenericC      74109 A74LS109DA2               DIP1674LS109D74LS109D                                                                  �    ����AA       ���������   ����AA      ���������   ����AA      ���������   ����AA      ��������InputInput                              �    ����AA     INA�  �  ClockClock                �    ����inIn     IN1A�  �>  �   ����outY     OUT1Y�  �>   �   &� 1 in   A1A&� 2 out   A1Y&� 3 in   B2A&� 4 out   B2Y&� 5 in   C3A&� 6 out   C3Y&� 7  GND  COMGND&� 8 out   D4Y&� 9 in  	 D4A&� 10 out  
 E5Y&� 11 in   E5A&� 12 out   F6Y&� 13 in   F6A&� 14  VCC  COMVCCdigital one-bit-wide inverterGatesGeneric=      7404 A74LS04DA3                                DIP1474LS04D74LS04D7�       inout 9� �>  in����    �  in����                         ��9� �>  out����   �  out����                        ��7404 LS Inverter7404 LS Inverter  8               }~Digital<   Generic                       * time value inInoutY IninYout                        �    ����AA     INA  Q  InputInput                  �    ����AA     INA  Q  InputInput                  �    ����portport       ��������Output_PortOutput_Port                  �    ����portport       ��������Output_PortOutput_Port                  �    ����portport       ��������Output_PortOutput_Port                �    ����SS     INS�      �   ����JJ     INJ�     �   ����ClkClk     INClk�     �   ����KK     INK�     �   ����RR     INR�     �   ����QQ     OUTQ�     �   ����Q'Q'     TRIQ'�      O �   WXYZ[\]^_`abcdef2JK pos edge triggered flip-flop w/preset and clear
Flip FlopsGenericC      74109 A74LS109DA2               DIP1674LS109D74LS109D                                                                  �    ����portport       ��������Output_PortOutput_Port                                                          p�t