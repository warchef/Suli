    � B2SPICE zzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzz 
 
 
 ��  CPart        �      p      �      p              74ALS192 (XSpice)��  CIntPin    ��  CWire       ��  	 TModelPin e
  Clr����        Clr����                          ��      x��    ��������      x��    ��������      x��    ��������      x��    ��������      x��    ��������      x��    �������� d   :�0�yE>10e-9��    �������� d   :�0�yE>10e-9��    ��������                             ����  ����:�0�yE>10e-9��d         ����  ����:�0�yE>10e-9��d   �      ��   T74192       ClrUpDownLoadABCDCOBOQAQBQCQD  � f
  Up����       Up����                          ��      x��    ��������      x��    ��������      x��    ��������      x��    ��������      x��    ��������      x��    �������� d   :�0�yE>10e-9��    �������� d   :�0�yE>10e-9��    ��������                            ����  ����:�0�yE>10e-9��d         ����  ����:�0�yE>10e-9��d   �     �    �       2    2
   �����     ��   d   :�0�yE>10e-9��    �������� d   :�0�yE>10e-9��    ��������� g
  Down����       Down����                          ��      x��    ��������      x��    ��������      x��    ��������      x��    ��������      x��    ��������      x��    �������� d   :�0�yE>10e-9��    �������� d   :�0�yE>10e-9��    ��������                            ����  ����:�0�yE>10e-9��d         ����  ����:�0�yE>10e-9��d   �     �    �       4 �        ��   TInPort       _   @         _   @                 Input ��  CExtPin    ��  CVertex   �  �	   ��  CSegment     �   `  �
                           @  �   A     `   	          In1     ��   CPin                    ��                                                       �   @   A��  TEllipse �   8   �   H                  ����
[negative]               ���                    �   8   �   H   �   8   �   H   �� 
 TRectangle t       �   @                   ����A                                      t       �   @   � t   @   �   `                   ����A                                      t   @   �   `   ��  TLine �   @   �   @     ��    ����                                                �         �   `                   ����                                                 �   `   "� t       t   `     
 ��    ����                                              ��  TPolygon                    ��                                                       ��  TPoint�   \        (��   P    �  (��   P    @  (��   D    ��S(��   D    �  (��   P    `  (��   P    P��    &�                    ��                                                       (��   $    `  (��   0    �  (��   0    �  (��   <       (��   <       (��   0       (��   0    ���    ��  
 TTextField �       �   8    	 ��        	                                               �       �   8   �       �   8   	[A.nbits]      <       ����            �      "Arial                �       �   8   8�    (      M     ��        
                                                 (      M      (      M   [value]       l  x	  �  
     (   l   P   8� ��������+   #     ��                                                       ��������+   #   ��������+   #   	[refname]       Z  �  �  �	  ���������        $   #   ! 0   : ' 9 ;      %      input_general     Miscellaneous      �?      ��   TInPortModel       A � Q  A����        A����                         ��             0��    ��������             0��    ��������             0��    ��������             0��    ��������             0��    ��������             0��    �������� d   :�0�yE>10e-9��    �������� d   :�0�yE>10e-9��    ��������                            ����  ����:�0�yE>10e-9��d         ����  ����:�0�yE>10e-9��d   �      =   �����        d   :�0�yE>10e-9��    �������� d   :�0�yE>10e-9��    ��������1 Bit Inport1 Bit Inport   �            > Digital<   Generic   In1In1           ����  ��    �������� ����  ��    �������� ����  ��    �������� ����  ��    �������� ����  ��    �������� ����  ��    �������� ����  ��    ��������  al      ����            In ��   CPartPin    ����AA      INAA�      Digital Instruments Generic                         `   `              `   �  �              `   �             �  `   `          �      4   >  4
   �����     ��   d   :�0�yE>10e-9��    �������� d   :�0�yE>10e-9��    ��������� h
  Load����       Load����                          ��      x��    ��������      x��    ��������      x��    ��������      x��    ��������      x��    ��������      x��    �������� d   :�0�yE>10e-9��    �������� d   :�0�yE>10e-9��    ��������                            ����  ����:�0�yE>10e-9��d         ����  ����:�0�yE>10e-9��d   �     �    �   B    5 �    B    �       _   @         _   @                 InputD �    �   `  �                    @  �   A        �
          In6     �                    ��                                                       �   @   A� �   8   �   H                  ����
[negative]               ���                    �   8   �   H   �   8   �   H   � t       �   @                   ����A                                      t       �   @   � t   @   �   `                   ����A                                      t   @   �   `   "� �   @   �   @     ��                                                        �         �   `                   ����                                                 �   `   "� t       t   `     
 ��                                                      &�                    ��                                                       (��   \        (��   P    �  (��   P    @  (��   D    ��S(��   D    �  (��   P    `  (��   P    P��    &�                    ��                                                       (��   $    `  (��   0    �  (��   0    �  (��   <       (��   <       (��   0       (��   0    ���    8� �       �   8    	 ��        	                                               �       �   8   �       �   8   	[A.nbits]      <       ����            �      "Arial                �       �   8   8�    (      M     ��        
                                                 (      M      (      M   [value]       ,  X  d  �     (   l   P   8� ��������+   #     ��                                                       ��������+   #   ��������+   #   	[refname]         �
  �  q  ���������       H M   L   K W   ` O _ a J   I N      input_general     Miscellaneous      �?      <�       A � Q  A����        A����                         ��             0��    ��������             0��    ��������             0��    ��������             0��    ��������             0��    ��������             0��    �������� d   :�0�yE>10e-9��    �������� d   :�0�yE>10e-9��    ��������                            ����  ����:�0�yE>10e-9��d         ����  ����:�0�yE>10e-9��d   �     B b   �����        d   :�0�yE>10e-9��    �������� d   :�0�yE>10e-9��    ��������1 Bit Inport1 Bit Inport   �            c Digital<   Generic   In6In6           ����  ��    �������� ����  ��    �������� ����  ��    �������� ����  ��    �������� ����  ��    �������� ����  ��    �������� ����  ��    ��������  ����    ����            In ?�    ����AA      INAA�?      Digital Instruments Generic               s G       `   `              `   �  �              `   �             �  `   `          �      5  A c  5
   �����     ��   d   :�0�yE>10e-9��    �������� d   :�0�yE>10e-9��    ��������� i
  A����       A����                          ��      x��    ��������      x��    ��������      x��    ��������      x��    ��������      x��    ��������      x��    �������� d   :�0�yE>10e-9��    �������� d   :�0�yE>10e-9��    ��������                             ����  ����:�0�yE>10e-9��d         ����  ����:�0�yE>10e-9��d   �     �    �   f    6 �    f    �       _   @         _   @                 Inputh �    �   �  `   �   k �   `  `   l                        @  �   A �a @  �          In2     �                    ��                                                       �   @   A� �   8   �   H                  ����
[negative]               ���                    �   8   �   H   �   8   �   H   � t       �   @                   ����A                                      t       �   @   � t   @   �   `                   ����A                                      t   @   �   `   "� �   @   �   @     ��                                                        �         �   `                   ����                                                 �   `   "� t       t   `     
 ��                                                      &�                    ��                                                       (��   \        (��   P    �  (��   P    @  (��   D    ��S(��   D    �  (��   P    `  (��   P    P��    &�                    ��                                                       (��   $    `  (��   0    �  (��   0    �  (��   <       (��   <       (��   0       (��   0    ���    8� �       �   8    	 ��        	                                               �       �   8   �       �   8   	[A.nbits]      <       ����            �      "Arial                �       �   8   8�    (      M     ��        
                                                 (      M      (      M   [value]       L    �  �     (   l   P   8� ��������+   #     ��                                                       ��������+   #   ��������+   #   	[refname]       :  �  �  1  ���������       n s   r   q }   � u � � p   o t      input_general     Miscellaneous      �?      <�       A � Q  A����        A����                         ��             0��    ��������             0��    ��������             0��    ��������             0��    ��������             0��    ��������             0��    �������� d   :�0�yE>10e-9��    �������� d   :�0�yE>10e-9��    ��������                            ����  ����:�0�yE>10e-9��d         ����  ����:�0�yE>10e-9��d   �     f �   �����         d   :�0�yE>10e-9��    �������� d   :�0�yE>10e-9��    ��������1 Bit Inport1 Bit Inport   �            � Digital<   Generic   In2In2           ����  ��    �������� ����  ��    �������� ����  ��    �������� ����  ��    �������� ����  ��    �������� ����  ��    �������� ����  ��    ��������          ����             In ?�    ����AA      INAA�?      Digital Instruments Generic                         `   `              `   �  �              `   �             �  `   `          �      6  e �  6
   �����     ��   d   :�0�yE>10e-9��    �������� d   :�0�yE>10e-9��    ��������� j
  B����       B����                          ��      x��    ��������      x��    ��������      x��    ��������      x��    ��������      x��    ��������      x��    �������� d   :�0�yE>10e-9��    �������� d   :�0�yE>10e-9��    ��������                             ����  ����:�0�yE>10e-9��d         ����  ����:�0�yE>10e-9��d   �     �    �   �    7 �    �    �       _   @         _   @                 Input� �    �   �      �   �   �  �   � �   � �   `  �   �                 �                @  �   A�Z�K @  `          In3     �                    ��                                                       �   @   A� �   8   �   H                  ����
[negative]               ���                    �   8   �   H   �   8   �   H   � t       �   @                   ����A                                      t       �   @   � t   @   �   `                   ����A                                      t   @   �   `   "� �   @   �   @     ��                                                        �         �   `                   ����                                                 �   `   "� t       t   `     
 ��                                                      &�                    ��                                                       (��   \        (��   P    �  (��   P    @  (��   D    ��S(��   D    �  (��   P    `  (��   P    P��    &�                    ��                                                       (��   $    `  (��   0    �  (��   0    �  (��   <       (��   <       (��   0       (��   0    ���    8� �       �   8    	 ��        	                                               �       �   8   �       �   8   	[A.nbits]      <       ����            �      "Arial                �       �   8   8�    (      M     ��        
                                                 (      M      (      M   [value]       L  �  �  n     (   l   P   8� ��������+   #     ��                                                       ��������+   #   ��������+   #   	[refname]       :  Q  �  �  ���������       � �   �   � �   � � � � �   � �      input_general     Miscellaneous      �?      <�       A � Q  A����        A����                         ��             0��    ��������             0��    ��������             0��    ��������             0��    ��������             0��    ��������             0��    �������� d   :�0�yE>10e-9��    �������� d   :�0�yE>10e-9��    ��������                            ����  ����:�0�yE>10e-9��d         ����  ����:�0�yE>10e-9��d   �     � �   �����         d   :�0�yE>10e-9��    �������� d   :�0�yE>10e-9��    ��������1 Bit Inport1 Bit Inport   �            � Digital<   Generic   In3In3           ����  ��    �������� ����  ��    �������� ����  ��    �������� ����  ��    �������� ����  ��    �������� ����  ��    �������� ����  ��    ��������          ����             In ?�    ����AA      INAA�?      Digital Instruments Generic                         `   `              `   �  �              `   �             �  `   `          �      7  � �  7
   �����     ��   d   :�0�yE>10e-9��    �������� d   :�0�yE>10e-9��    ��������� k
  C����       C����                          ��      x��    ��������      x��    ��������      x��    ��������      x��    ��������      x��    ��������      x��    �������� d   :�0�yE>10e-9��    �������� d   :�0�yE>10e-9��    ��������                             ����  ����:�0�yE>10e-9��d         ����  ����:�0�yE>10e-9��d   �     �    �   �    8 �    �    �       _   @         _   @                 Input� �    �   �  �   �   � �   �  �   � �   �   �      � �   � �   `      �                 �                        @  �   A �a @             In4     �                    ��                                                       �   @   A� �   8   �   H                  ����
[negative]               ���                    �   8   �   H   �   8   �   H   � t       �   @                   ����A                                      t       �   @   � t   @   �   `                   ����A                                      t   @   �   `   "� �   @   �   @     ��                                                        �         �   `                   ����                                                 �   `   "� t       t   `     
 ��                                                      &�                    ��                                                       (��   \        (��   P    �  (��   P    @  (��   D    ��S(��   D    �  (��   P    `  (��   P    P��    &�                    ��                                                       (��   $    `  (��   0    �  (��   0    �  (��   <       (��   <       (��   0       (��   0    ���    8� �       �   8    	 ��        	                                               �       �   8   �       �   8   	[A.nbits]      <       ����            �      "Arial                �       �   8   8�    (      M     ��        
                                                 (      M      (      M   [value]       L  �  �  .     (   l   P   8� ��������+   #     ��                                                       ��������+   #   ��������+   #   	[refname]       :    �  �  ���������       � �   �   � �   � � � � �   � �      input_general     Miscellaneous      �?      <�       A � Q  A����        A����                         ��             0��    ��������             0��    ��������             0��    ��������             0��    ��������             0��    ��������             0��    �������� d   :�0�yE>10e-9��    �������� d   :�0�yE>10e-9��    ��������                            ����  ����:�0�yE>10e-9��d         ����  ����:�0�yE>10e-9��d   �     � �   �����         d   :�0�yE>10e-9��    �������� d   :�0�yE>10e-9��    ��������1 Bit Inport1 Bit Inport   �            � Digital<   Generic   In4In4           ����  ��    �������� ����  ��    �������� ����  ��    �������� ����  ��    �������� ����  ��    �������� ����  ��    �������� ����  ��    ��������         ����             In ?�    ����AA      INAA�?      Digital Instruments Generic                         `   `              `   �  �              `   �             �  `   `          �      8  � �  8
   �����     ��   d   :�0�yE>10e-9��    �������� d   :�0�yE>10e-9��    ��������� l
  D����       D����                          ��      x��    ��������      x��    ��������      x��    ��������      x��    ��������      x��    ��������      x��    �������� d   :�0�yE>10e-9��    �������� d   :�0�yE>10e-9��    ��������                             ����  ����:�0�yE>10e-9��d         ����  ����:�0�yE>10e-9��d   �     �    �   �    9 �    �    �       _   @         _   @                 Input� �    �   �  �   �   � �   `  �   � �   �   `  �   �         �                        @  �   AY�K @  �          In5     �                    ��                                                       �   @   A� �   8   �   H                  ����
[negative]               ���                    �   8   �   H   �   8   �   H   � t       �   @                   ����A                                      t       �   @   � t   @   �   `                   ����A                                      t   @   �   `   "� �   @   �   @     ��                                                        �         �   `                   ����                                                 �   `   "� t       t   `     
 ��                                                      &�                    ��                                                       (��   \        (��   P    �  (��   P    @  (��   D    ��S(��   D    �  (��   P    `  (��   P    P��    &�                    ��                                                       (��   $    `  (��   0    �  (��   0    �  (��   <       (��   <       (��   0       (��   0    ���    8� �       �   8    	 ��        	                                               �       �   8   �       �   8   	[A.nbits]      <       ����            �      "Arial                �       �   8   8�    (      M     ��        
                                                 (      M      (      M   [value]       L  X  �  �     (   l   P   8� ��������+   #     ��                                                       ��������+   #   ��������+   #   	[refname]       :  �  �  q  ���������       � �   �   � �    � � �   � �      input_general     Miscellaneous      �?      <�       A � Q  A����        A����                         ��             0��    ��������             0��    ��������             0��    ��������             0��    ��������             0��    ��������             0��    �������� d   :�0�yE>10e-9��    �������� d   :�0�yE>10e-9��    ��������                            ����  ����:�0�yE>10e-9��d         ����  ����:�0�yE>10e-9��d   �     �   �����         d   :�0�yE>10e-9��    �������� d   :�0�yE>10e-9��    ��������1 Bit Inport1 Bit Inport   �            Digital<   Generic   In5In5           ����  ��    �������� ����  ��    �������� ����  ��    �������� ����  ��    �������� ����  ��    �������� ����  ��    �������� ����  ��    ��������         ����             In ?�    ����AA      INAA�?      Digital Instruments Generic               0��       `   `              `   �  �              `   �             �  `   `          �      9  �  9
   �����     ��   d   :�0�yE>10e-9��    �������� d   :�0�yE>10e-9��    ��������� m
  CO����       CO����                         �� �   h�+e�SS>18ns��    �������� 2   :�0�y5>5ns��    ��������      x��    �������� �   ��&�.Q>16ns��    �������� (   ��&�.1>4ns��    ��������      x��    �������� d   :�0�yE>10e-9��    �������� d   :�0�yE>10e-9��    ��������                           ����  ����:�0�yE>10e-9��d         ����  ����:�0�yE>10e-9��d   �     �    �      10   10
   �����          d   :�0�yE>10e-9��    �������� d   :�0�yE>10e-9��    ��������� n
  BO����	       BO����                         �� �   h�+e�SS>18ns��    �������� 2   :�0�y5>5ns��    ��������      x��    �������� �   ,i�)+P>15ns��    �������� (   ��&�.1>4ns��    ��������      x��    �������� d   :�0�yE>10e-9��    �������� d   :�0�yE>10e-9��    ��������                           ����  ����:�0�yE>10e-9��d         ����  ����:�0�yE>10e-9��d   �     �	    �	   		 	  11  	 11
   �����          d   :�0�yE>10e-9��    �������� d   :�0�yE>10e-9��    ��������� o
  QA����
       QA����                         ��   ��C֔^>28ns��    �������� 9   �$^7{8>5.7ns��    ��������      x��    �������� ,  ,i�)+`>30ns��    �������� <   �A:��9>6ns��    ��������      x��    �������� d   :�0�yE>10e-9��    �������� d   :�0�yE>10e-9��    ��������                            ����  ����:�0�yE>10e-9��d         ����  ����:�0�yE>10e-9��d   �     �
    �
   
 
  12  
 12
   �����     ��  d   :�0�yE>10e-9��    �������� d   :�0�yE>10e-9��    ��������� p
  QB����       QB����                         ��   ��C֔^>28ns��    �������� 9   �$^7{8>5.7ns��    ��������      x��    �������� ,  ,i�)+`>30ns��    �������� <   �A:��9>6ns��    ��������      x��    �������� d   :�0�yE>10e-9��    �������� d   :�0�yE>10e-9��    ��������                            ����  ����:�0�yE>10e-9��d         ����  ����:�0�yE>10e-9��d   �     �    �      13 �      �       �   �  p      �   �  p              74LS08N�   �    �      15  � r
  QD����       QD����                         ��   ��C֔^>28ns��    �������� 9   �$^7{8>5.7ns��    ��������      x��    �������� ,  ,i�)+`>30ns��    �������� <   �A:��9>6ns��    ��������      x��    �������� d   :�0�yE>10e-9��    �������� d   :�0�yE>10e-9��    ��������                            ����  ����:�0�yE>10e-9��d         ����  ����:�0�yE>10e-9��d   �     
   �����     ��  d   :�0�yE>10e-9��    �������� d   :�0�yE>10e-9��    ��������� <  B����       B����                          ��      x��    ��������      x��    ��������      x��    ��������      x��    ��������      x��    ��������      x��    �������� d   :�0�yE>10e-9��    �������� d   :�0�yE>10e-9��    ��������                             ����  ����:�0�yE>10e-9��d         ����  ����:�0�yE>10e-9��d   �     ��   TAnd       ABY � ;  A����        A����                          ��      x��    ��������      x��    ��������      x��    ��������      x��    ��������      x��    ��������      x��    �������� d   :�0�yE>10e-9��    �������� d   :�0�yE>10e-9��    ��������                             ����  ����:�0�yE>10e-9��d         ����  ����:�0�yE>10e-9��d   �       �����     ��   d   :�0�yE>10e-9��    �������� d   :�0�yE>10e-9��    ��������� =  Y����       Y����                         �� �   :�0�yU>20ns��    ��������      x��    �������� d   :�0�yE>10ns��    �������� �   ,i�)+P>15ns��    ��������      x��    �������� P   ��&�.A>8ns��    �������� d   :�0�yE>10e-9��    �������� d   :�0�yE>10e-9��    ��������                            ����  ����:�0�yE>10e-9��d         ����  ����:�0�yE>10e-9��d   �     �    �      16 �       ��   TOutPort	       _   @         _   @                 Output_Port�    �   �               	            �   port     �  `          Out2     �                   ��                                                           @   port�         �   `                   ����                                                 �   `   "�     @       @      ��                                                        �    8       H                  ����
[negative]               ���                       8       H      8       H   8� (   ,   E   Q     ��                                                      (   ,   E   Q   (   ,   E   Q   [value]       X  �  �  z  (   ,   �   T   8�     $       <     ��                                                           $       <       $       <   [port.nbits]      <       ����            �      "Arial                    $       <   8�     ����j         ��                                                           ����j           ����j       	[refname]       @  H     �      �����       %  #&'()$     Output_Port     Miscellaneous      �?      ��   TOutPortModel       port � ����port����        port����                                         0��    ��������             0��    ��������             0��    ��������             0��    ��������             0��    ��������             0��    �������� d   :�0�yE>10e-9��    �������� d   :�0�yE>10e-9��    ��������                             ����  ����:�0�yE>10e-9��d         ����  ����:�0�yE>10e-9��d   �     +  �����     ��   d   :�0�yE>10e-9��    �������� d   :�0�yE>10e-9��    ��������Output_PortOutput_Port   �            ,Digital<   Generic   Out2Out2           ����  ��    �������� ����  ��    �������� ����  ��    �������� ����  ��    �������� ����  ��    �������� ����  ��    �������� ����  ��    ��������  ���t    ����       ����  Out ?�    ����portport       A �?      Digital Instruments Generic                                                                          yE>                                16  , 16  �����     ��  d   :�0�yE>10e-9��    �������� d   :�0�yE>10e-9��    ��������08/4 LS 2-Inp. And08/4 LS 2-Inp. And  A �t            Digital<   Analog Devices   A2A2           ���� x��    �������� ���� x��    �������� @ �h㈵��>20u��    �������� ���-C��6:�-.4m��    �������� ���-C��6:�-.4m��    ��������  ������Mb�?8m��    �������� ��`�Q�k?3.4m��    ��������  ��&�    ����LS      �����     ��   d   :�0�yE>10e-9��    �������� d   :�0�yE>10e-9��    �������� 15  15 �    "  �  �  y    �   �      �   �	   �   �
  �   1        0    �
   0�   `  �   3                         a   �   �      �   �   �   �
  �   �   �    
  �   9    8    7        6                 �  b       �          A2     �                   ��                                                       �   �   y�                    ��                                                          `   a�                   ��                                                          �   b"�     P       �    
 ��                                                        "�     �       �    	 ��                                                        "�     `       `     ��                                                        "� �   �   �   �     ��                                                        "�     �   D   �     ��    ����                                                ��   TArc    P   �   �                                                                  P   �   �      P   �   �   �   �   D   P           "�     P   D   P     ��    ����	                                                C�    0   �   �               
                                                   0   �   �      0   �   �   D   �   �   �           8�     �����        ��                                                           �����          �����      	[devname]        ����������������    �����      8�        b   D     ��                                                              b   D          b   D   	[refname]       `  �  (  �         �   @    <=  F  E;D  B  HAG  @  ?  >     AND 2    
AND 2 IEEEMiscellaneous      �?    A    A ?�    ����aA      INA1A����    ?�   ����bB      INA1B�?     ?�   ����yY      OUTA1Y8@     ?�    ����aA      INB1A7@      ?�   ����bB      INB1B6@     ?�   ����yY      OUTB1Y�?     ?�    ����aA      INC1A�?      ?�   ����bB      INC1B�?     ?�   ����yY      OUTC1Y       ?�    ����aA      IND1A�?      ?�   ����bB      IND1B�?     ?�   ����yY      OUTD1Y�>     GatesXSpice 2input AND gateGenericDIP-14              13   13
   �����     ��  d   :�0�yE>10e-9��    �������� d   :�0�yE>10e-9��    ��������� q
  QC����       QC����                         ��   ��C֔^>28ns��    �������� 9   �$^7{8>5.7ns��    ��������      x��    �������� ,  ,i�)+`>30ns��    �������� <   �A:��9>6ns��    ��������      x��    �������� d   :�0�yE>10e-9��    �������� d   :�0�yE>10e-9��    ��������                            ����  ����:�0�yE>10e-9��d         ����  ����:�0�yE>10e-9��d   �     �    �   V   14  U 14
   �����     ��  d   :�0�yE>10e-9��    �������� d   :�0�yE>10e-9��    ��������192 ALS Up/Down Counter192 ALS Up/Down Counter  b T               A e � � � UDigital<   Motorola   A1A1           ���� x��    �������� ���� x��    �������� @ �h㈵��>20u��    �������� �{��-C��6*�-.2m��    �������� ���-C��6:�-.4m��    ��������  ������Mb�?8m��    ��������  '�~j�t��?12m��    ��������  V l     ����ALS        �A:��>1.5n��    �������� ����    ��wA25meg��    �������� �   �C���@R>17n��    �������� �   :�0�yU>20n��    ��������  �����     ��   d   :�0�yE>10e-9��    �������� d   :�0�yE>10e-9��    ��������  3  �� 3   C g � � � 
W�    �    `  �	                     �  Clr    �   �   `   
                  �  Up   �          �  Down   �   G       `  Load   �   m          A   �   �       �  B   �   �       �  C   �   �       @  D   �   �   �
   
                 �  CO   �	   �	   �
  �
     	      	  	    �  BO	   �
   �
   �
  `     
      
  
       QA
   �   2     �  QB   �   �   �
                    �  QC   �   8     @  QD    `  @          A1    A �                   ��                                                           �   Clr�                   ��                                                          �   Up�                   ��                                                          �   Down�                   ��                                                             Load�                   ��                                                          `  A�                   ��                                                          �  B�                   ��                                                          �  C�                   ��                                                          �  D�                  	 ��                                                      `  �   CO�                  
 ��        	                                              `  �   BO�                   ��        
                                              `  `  QA�                   ��                                                      `  �  QB�                   ��                                                      `  �  QC�                   ��                                                      `  �  QD� @   P     �                 ����                                         @   P     �  "�     �   @   �     ��       �                                                "�     �   @   �     ��     	                                                  "�     �   @   �     ��    `	                                                  "�    �   4  �    . ��                                                        "�    �      �    / ��    8�b                                                "�     �           3 ��    �	                                                  "�        @       2 ��    	                                                   "�     �   @   �    1 ��    �� �                                                "�     �       �    0 ��    �                                                  "� @   p     p   6 ��                                                       "� @   �     �   7 ��                                                        "� @   �     �   8 ��                                                        "� �   �   �   �    = ��                                                        "� �   �   �   �    > ��                                                        "�        @        ��                                                        "�     `  @   `    ��    ��W                                                "�     �  @   �    ��                                                        "�     �  @   �    ��    H                                                   "�     �  @   �    ��    X�R!                                                "�    �   `  �     ��    \  "                                                "�    �   `  �     ��    p�R#                                                "�    `  `  `    ��    �� �$                                                "�    �  `  �    ��    4�R%                                                "�    �  `  �    ��    ��[&                                                "�    �  `  �    ��    �,b'                                                "� @   �   L   �    & ��    (Y](                                                "� L   �   @   �    ' ��    �  )                                                "� L   �   @   �    ( ��    �Y*                                                "� @   �   L   �    ) ��    �  +                                                "� ,     ,       * ��    Z],                                                "� ,     @       + ��    �  -                                                "�    �   4  �    , ��    X.b.                                                "�    �      �    - ��    �  /                                                &� ����������������   ��        0                                                 (�P   P  0  2[(�P   @  0     (�@   @  0     (�@   @   0     (�   @   0     (�   @  0     (�  @  0 �T(�  P  0         8� H   p   �   �     ��        1                                              H   p   �   �   H   p   �   �   ct=0       8  �	  �  &
  H   p   �   �   8� T   �   y   �     ��        2                                              T   �   y   �   T   �   y   �   2+       \  �	  �  �
  T   �   |   �   8� T   �   q   �      ��        3                                              T   �   q   �   T   �   q   �   1-       \  �
  �  F  T   �   |   �   8� H     j   5   ! ��        4                                              H     j   5  H     j   5  c3       8  p  �    H     �   0  8� H   P  m   u   " ��        5                                              H   P  m   u  H   P  m   u  3d       8  0  �  �  H   P  t   p  8� h   @   �   e    # ��        6                                              h   @   �   e   h   @   �   e   	ctrdIv 10       �   	   	  �	  h   @     `   8� H   �   m   �    4 ��        7                                              H   �   m   �   H   �   m   �   g1       8  P
  �  �
  H   �   p   �   8� �   �     �    $ ��        8                                              �   �     �   �   �     �   1ct=9       �  �	  �	  �
  �   �      �   8� �   �     �    % ��        9                                              �   �     �   �   �     �   2ct=0       �  �
  �	  F  �   �      �   8� H   �   m      5 ��        :                                              H   �   m     H   �   m     g2       8    �  �  H   �   p     8� �   L  �   q   9 ��        ;                                              �   L  �   q  �   L  �   q  [1]       L  $  �  �  �   L  �   l  8� �   l  �   �   : ��        <                                              �   l  �   �  �   l  �   �  [2]       L  �  �    �   l  �   �  8� �   �  �   �   ; ��        =                                              �   �  �   �  �   �  �   �  [4]       L  �  �  z  �   �  �   �  8� �   �  �   �   < ��        >                                              �   �  �   �  �   �  �   �  [8]       L  D  �  �  �   �  �   �  8� @      j   <    ? ��        ?                                               @      j   <   @      j   <   	[refname]          |  �  	  @      �   8   8� @   �����       @ ��        @                                               @   �����      @   �����      	[devname]        ����������������@   �����      c �  lmnopqrstuvwxyz{|}�������������������                ��������������    ��                                  ~�  �  �  ����      ���     74192 Up/Down Counter     Miscellaneous      �?    b  
   A ?�    ����ClrClr      INAClr        ?�   ����UpUp      INAUp       ?�   ����DownDown      INADownӑ)A   ?�   ����LoadLoad      INALoad> �r   ?�   ����AA      INAAB�r   ?�   ����BB      INAB       ?�   ����CC      INAC����   ?�   ����DD      INAD�� �   ?�   ����COCO      OUTACO      ?�	   ����BOBO      OUTABO    	   ?�
   ����QAQA      OUTAQA    
   ?�   ����QBQB      OUTAQB��Y	   ?�   ����QCQC      OUTAQC       ?�   ����QDQD      OUTAQD       Counters(synchronous 4-bit up/down decade counterGeneric                i � � � E �       _   @         _   @                   Output_Port�    �   `�                       �   port     `�  `          Out1     �                   ��                                                           @   port�         �   `                   ����                                                 �   `   "�     @       @      ��                                                        �    8       H                  ����
[negative]               ���                       8       H      8       H   8� (   ,   �   T     ��                                                      (   ,   `   Q   (   ,   `   Q   [value]       ��  �  ��  z  (   ,   �   T   8�     $       <     ��                                                           $       <       $       <   [port.nbits]      <       ����            �      "Arial                    $       <   8�     �����        ��                                                           ����j           ����j       	[refname]       ��  H  ��  �      �����       �  ������     Output_Port     Miscellaneous      �?      *�       port  Output_PortOutput_Port   �             Digital<   Generic   Out1Out1           ����  ��    �������� ����  ��    �������� ����  ��    �������� ����  ��    �������� ����  ��    �������� ����  ��    �������� ����  ��    ��������  d       ����       ����  Out  Digital Instruments Generic                                                                                                                    B f � � � 	V    l � � � � � � � 1397         Y[k G � � � � ceg2j8  � � m � � � � "06�4:                 
 ��  CValue@ ����        ��������΁             0     ��������΁ ����      @5     ��������΁  ʚ;�������?.1     ��������΁@ ����       ��������΁ ����       ��������΁ ����       ��������΁ ����       ��������΁ ���� true
     ��������΁ ����  false     ��������               
                  ΁ ����        ��������΁ ����       ��������΁  ����       ��������΁@ ����       ��������΁@ ����       ��������               
                  ΁ ����        ��������΁ ����       ��������΁@ ����       ��������΁  ����       ��������΁ ����       ��������΁ ����       ��������΁ ����       ��������΁ ����       ��������΁ ����       ��������΁ ����       ��������΁ ����       ��������               
                 ΁ ����dec     ��������΁ ����     @�@1k     ��������΁ ����    ��.A1meg     ��������΁ ����       20     ��������΁ ���� true     ��������΁ ���� true     ��������΁ ���� true	     ��������΁ ����  false
     ��������               
                 ΁  ����        ��������΁  ����       ��������΁  ����       ��������΁ ����dec     ��������΁ ����       ��������΁ ����       ��������΁ ����  	     ��������΁ ����  
     ��������               
                  	 ΁ ����        ��������΁ ����       ��������΁ ����       ��������΁ ����       ��������΁ ����       ��������΁ ����       ��������΁ ����       ��������΁ ����       ��������΁ ����       ��������               
                 ΁ ����        ��������΁ ����       ��������΁ ����       ��������΁ ����dec     ��������΁ ����       ��������               
                    ΁             0      ��������΁ ��� ����MbP?1m     ��������΁ �� �h㈵��>10u     ��������΁ '  ���ư>1u     ��������΁ ���� true     ��������΁ ����  false     ��������΁ ���� true     ��������΁ ����  false     ��������               
                 ΁ ����     @�@1K      ��������΁  ����       ��������΁  ����       ��������΁  ����       ��������               
         ��              ΁  ����        ��������              
                  ΁  ����        ��������              
                                  
                 ΁@ ����        ��������΁@ ����       ��������΁ ����       ��������΁ ����       ��������΁ ����       ��������΁ ����       ��������΁ ����       ��������΁ ����       ��������΁ ����       ��������΁ ���� true	     ��������΁ ����  false
     ��������΁ ���� true     ��������΁ ����  false     ��������               
                 ΁ ����       5      ��������΁ ����       5     ��������΁ ����       5     ��������΁ ����       5     ��������΁ ����       ��������΁ ����  	     ��������΁ ����  
     ��������΁ ����       ��������΁ ����       ��������΁ ����       ��������΁ ���� true     ��������΁@ ����       ��������΁@ ����       ��������΁ ����       ��������΁ ����       ��������΁ ����       ��������΁ ����dec     ��������΁ ����       ��������΁ ����       ��������΁ ����       ��������΁ ���� true     ��������΁ ���� true     ��������΁ ���� true     ��������΁ ����  false     ��������΁ ���� true     ��������΁ ����  false      ��������΁ ���� true!     ��������΁ ����  false"     ��������               
                        ΁ ����       5      ��������΁ ����       5     ��������΁ ����       5     ��������΁ ����       5     ��������΁ ����       ��������΁ ����  	     ��������΁ ����  
     ��������΁ ����       ��������΁ ����       ��������΁ ����       ��������΁ ���� true     ��������΁@ ����       ��������΁@ ����       ��������΁ ����       ��������΁ ����       ��������΁ ����       ��������΁ ����dec     ��������΁ ����       ��������΁ ����       ��������΁ ����       ��������΁ ���� true     ��������΁ ���� true     ��������΁ ���� true     ��������΁ ����  false     ��������΁ ���� true     ��������΁ ����  false      ��������΁ ���� true!     ��������΁ ����  false"     ��������               
                 ΁ ����       5      ��������΁ ����       5     ��������΁ ����       5     ��������΁ ����       5     ��������΁ ����       ��������΁ ����  	     ��������΁ ����  
     ��������΁ ����       ��������΁ ����       ��������΁ ����       ��������΁ ���� true     ��������΁@ ����       ��������΁@ ����       ��������΁ ����       ��������΁ ����       ��������΁ ����       ��������΁ ����dec     ��������΁ ����       ��������΁ ����       ��������΁ ����       ��������΁ ���� true     ��������΁ ���� true     ��������΁ ���� true     ��������΁ ����  false     ��������΁ ���� true     ��������΁ ����  false      ��������΁ ���� true!     ��������΁ ����  false"     ��������               
                 ΁ ����       5      ��������΁ ����       5     ��������΁ ����       5     ��������΁ ����       5     ��������΁ ����       ��������΁ ����  	     ��������΁ ����  
     ��������΁ ����       ��������΁ ����       ��������΁ ����       ��������΁ ���� true     ��������΁@ ����       ��������΁@ ����       ��������΁ ����       ��������΁ ����       ��������΁ ����       ��������΁ ����dec     ��������΁ ����       ��������΁ ����       ��������΁ ����       ��������΁ ���� true     ��������΁ ���� true     ��������΁ ���� true     ��������΁ ����  false     ��������΁ ���� true     ��������΁ ����  false      ��������΁ ���� true!     ��������΁ ����  false"     ��������               
                 ΁@ ����        ��������΁@ ����       ��������΁ ����       ��������΁ ����       ��������΁ ����       ��������΁ ����       ��������΁ ����       ��������΁ ����       ��������΁ ����decade     ��������΁ ���� true     ��������΁ ���� true     ��������΁ ���� true     ��������΁ ����  false     ��������               
                 ΁ ����        ��������΁ ����       ��������΁@ ����       ��������΁  ����       ��������΁ ����       ��������΁ ����       ��������΁ ����       ��������΁ ����       ��������΁ ����       ��������΁ ����       ��������΁ ����       ��������               
                        ΁ ����dec     ��������΁ ����     @�@1k     ��������΁ ����    ��.A1meg     ��������΁ ����       20     ��������΁ ����        0     ��������΁ ����        0     ��������΁ ���� true	     ��������΁ ���� true
     ��������΁ ����      I@50     ��������΁ ���� true     ��������΁ ����  false     ��������               
                          / ΁ ���� x'     ��������΁     �-���q=1E-12     ��������΁ @B -C��6?1E-4     ��������΁ ���� x     ��������΁ ���� x     ��������΁ ���� x     ��������΁ ���� x     ��������΁ ���� x     ��������΁ ���� x     ��������΁ ���� x	     ��������΁ ���� x!     ��������΁ ����    �  500
     ��������΁ ���� x     ��������΁ ����    �  500     ��������΁ ���� x$     ��������΁ ���� x$     ��������΁ ���� x%     ��������΁ ���� x"     ��������΁  ���� x*     ��������΁ ���� x     ��������΁ ���� x     ��������΁ ���� x     ��������΁ ���� x&     ��������΁ ���� x     ��������΁ ���� x     ��������΁ ���� x     ��������΁ ���� x+     ��������΁ ���� x,     ��������΁ ���� x-     ��������΁ ���� xg     ��������΁ ���� xf     ��������΁ ���� xd     ��������΁ ���� xe     ��������΁ ���� xh     ��������΁ ���� xj     ��������΁ ���� xi     ��������΁ ���� xk     ��������΁ ����    e��A1Gl     ��������΁             0�     ��������΁ ����      @5�     ��������΁ ����      @2.5�     ��������΁ ����      �?.5�     ��������΁ ����      @4.5�     ��������΁ 
   ��&�.>1n�     ��������΁ 
   ��&�.>1n�     ��������΁ 
   ��&�.>1n�     ��������΁ 
   ��&�.>1n�     ��������                                  Ariald        �ڬt4�e|�  ۬t0� ���t    �ڬt4�e|�  ۬t0� ���t ��  COpAnal                         
                        ����            `j�                   �ڬt4�e|�  ۬t0� ���t    �ڬt4�e|�  ۬t0� ���t ��  CDCsweep       
 ����������               
                      ����            ����                   �ڬt4�e|�  ۬t0� ���t    �ڬt4�e|�  ۬t0� ���t ��  CACsweep        ��������               
                      ����           �g�                   �ڬt4�e|�  ۬t0� ���t    �ڬt4�e|�  ۬t0� ���t �� 
 CTranSweep        	
               
                      ����            �  �                   �ڬt4�e|�  ۬t0� ���t    �ڬt4�e|�  ۬t0� ���t ��  CACdisto                       
                         ����                                 �ڬt4�e|�  ۬t0� ���t    �ڬt4�e|�  ۬t0� ���t �        ΁ ����        ��������΁ ����       ��������΁ ����       ��������΁ ����dec     ��������΁ ����       ��������               
                         ����            �v                    �ڬt4�e|�  ۬t0� ���t    �ڬt4�e|�  ۬t0� ���t �        ΁ ����        ��������΁ ����       ��������΁ ����       ��������΁ ����dec     ��������΁ ����       ��������               
                         ����                                 �ڬt4�e|�  ۬t0� ���t    �ڬt4�e|�  ۬t0� ���t �        ΁ ����        ��������΁ ����       ��������΁ ����       ��������΁ ����dec     ��������΁ ����       ��������               
                         ����                                  �ڬt4�e|�  ۬t0� ���t    �ڬt4�e|�  ۬t0� ���t �        ΁ ����        ��������΁ ����       ��������΁ ����       ��������΁ ����dec     ��������΁ ����       ��������               
                          ����                                 �ڬt4�e|�  ۬t0� ���t    �ڬt4�e|�  ۬t0� ���t �        ΁ ����        ��������΁ ����       ��������΁ ����       ��������΁ ����dec     ��������΁ ����       ��������               
         �            	    ����             ��                   �ڬt4�e|�  ۬t0� ���t    �ڬt4�e|�  ۬t0� ���t ��  CACnoise        ��������               
                   
    ����                                  �ڬt4�e|�  ۬t0� ���t    �ڬt4�e|�  ۬t0� ���t �                        
                        ����                                  �ڬt4�e|�  ۬t0� ���t    �ڬt4�e|�  ۬t0� ���t ��  CFourier                       
         ��                  ����                                  �ڬt4�e|�  ۬t0� ���t    �ڬt4�e|�  ۬t0� ���t ��  CACpz        	 �������                
                       ����                                   �ڬt4�e|�  ۬t0� ���t    �ڬt4�e|�  ۬t0� ���t ��  CDCtf         �����               
                       ����             x�                   �ڬt4�e|�  ۬t0� ���t    �ڬt4�e|�  ۬t0� ���t ��  CDCsens         �����������               
                       ����            �� �                   �ڬt4�e|�  ۬t0� ���t    �ڬt4�e|�  ۬t0� ���t                 ����            :                      �ڬt4�e|�  ۬t0� ���t    �ڬt4�e|�  ۬t0� ���t ��  CShow                       
                       ����            x� �                   �ڬt4�e|�  ۬t0� ���t    �ڬt4�e|�  ۬t0� ���t ��  CShowmod                       
                       ����            x��                   �ڬt4�e|�  ۬t0� ���t    �ڬt4�e|�  ۬t0� ���t �� 
 CLinearize        ΁  ����        ��������               
                      ����            �                     �ڬt4�e|�  ۬t0� ���t    �ڬt4�e|�  ۬t0� ���t ��  CParamTranSweep         !               
                      ����            �                     �ڬt4�e|�  ۬t0� ���t    �ڬt4�e|�  ۬t0� ���t �             ����                                  �ڬt4�e|�  ۬t0� ���t    �ڬt4�e|�  ۬t0� ���t ��  CParamACSweep        �������������               
                      ����           F                      �ڬt4�e|�  ۬t0� ���t    �ڬt4�e|�  ۬t0� ���t ��  CMonteCarlo_op        "#$%&'()*+,-./0123456789:;<=               
                             ����               �                   �ڬt4�e|�  ۬t0� ���t    �ڬt4�e|�  ۬t0� ���t ��  CMonteCarlo_dc        >?@ABCDEFGHIJKLMNOPQRSTUVWXY               
                      ����            x��                   �ڬt4�e|�  ۬t0� ���t    �ڬt4�e|�  ۬t0� ���t ��  CMonteCarlo_ac        Z[\]^_`abcdefghijklmnopqrstu               
                      ����           �                     �ڬt4�e|�  ۬t0� ���t    �ڬt4�e|�  ۬t0� ���t ��  CMonteCarlo_tran        vwxyz{|}~������������������               
                      ����                                  �ڬt4�e|�  ۬t0� ���t    �ڬt4�e|�  ۬t0� ���t ��  CACsens        �����������               
                             ����              �                   �ڬt4�e|�  ۬t0� ���t    �ڬt4�e|�  ۬t0� ���t ��  CNetworkAnalysis        �����������               
                      ����           x��                   �ڬt4�e|�  ۬t0� ���t    �ڬt4�e|�  ۬t0� ���t                 ����            �                   >           ��   CDigSimResTemplate                     ��   TDigitalSignal            In1    ���� ����                        0�            In2    ���� ����                        0�            In3    ���� ����                        0�            In4    ���� ����                        0�            In5    ���� ����                        0�            In6    ���� ����                        0�            Out1    ���� ����                         0�            Out2    ���� ����                              ��W���       ����  ����:�0�yU>+20.00n���   ����                       Arial����                       Arial����                       Arial                                           ����  ���� ������       ����  ���� ������                 �               ����  �����       200������          0.000000e+000��    ��������      0.000000e+000��    ��������      0.000000e+000��    ��������   ����                       Arial����                       Arial����                       Arial����                       Arial                        �     �   �  �                     ����  ��    ��������                                                                                                                 �   DIP-14�14 pin dual in line package                                                                                                                                                                                                                               �     ��   CPackageAliasSuperPCBStandardDIP14      9�EagleBURR.LBRDIP-14      9�Orcad DIP.100/14/W.300/L.700      9�Pads DIP14      9�	UltiboardUltilib.l55DIP14      9�Eagleburr-brown.lbrDIL14      9�Eagledil.lbrDIL14     9�Eagleanalog-devicesDIL14      9�Eagle74xx-usDIL14      9�Eagle	74ttl-dinDIL14      9�EaglemaximDIL14      9�EagleexarDIL14      9�Eagle
ic-packageDIL14      9�Eagleresistor-dilDIL14      9�EagletexasDIL14      9�Eagle
74ac-logicDIL14              A                            �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                   �#     ����x� H�]	    @�     J   J   ��     H�]	J                  2         �                 � � �           u m     ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                   �#     ����x� H�]	    @�     J   J   ��     H�]	J                  2         �                 � � �           u m     ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                   �#     ����x� H�]	    @�     J   J   ��     H�]	J                  2         �                 � � �           u m     ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                   �#     ����x� H�]	    @�     J   J   ��     H�]	J                  2         �                 � � �           u m     ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                   �#     ����x� H�]	    @�     J   J   ��     H�]	J                  2         �                 � � �           u m     ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                   �#     ����x� H�]	    @�     J   J   ��     H�]	J                  2         �                 � � �           u m     ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                   �#     ����x� H�]	    @�     J   J   ��     H�]	J                  2         �                 � � �           u m     ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                   �#     ����x� H�]	    @�     J   J   ��     H�]	J                  2         �                 � � �           u m     ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                   �#     ����x� H�]	    @�     J   J   ��     H�]	J                  2         �                 � � �           u m     ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                   �#     ����x� H�]	    @�     J   J   ��     H�]	J                  2         �                 � � �           u m     ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                   �#     ����x� H�]	    @�     J   J   ��     H�]	J                  2         �                 � � �           u m     ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                   �#     ����x� H�]	    @�     J   J   ��     H�]	J                  2         �                 � � �           u m     ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                   �#     ����x� H�]	    @�     J   J   ��     H�]	J                  2         �                 � � �           u m     ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                   �#     ����x� H�]	    @�     J   J   ��     H�]	J                  2         �                 � � �           u m     ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                   �#     ����x� H�]	    @�     J   J   ��     H�]	J                  2         �                 � � �           u m     ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                   �#     ����x� H�]	    @�     J   J   ��     H�]	J                  2         �                 � � �           u m     ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                   �#     ����x� H�]	    @�     J   J   ��     H�]	J                  2         �                 � � �           u m     ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                   �#     ����x� H�]	    @�     J   J   ��     H�]	J                  2         �                 � � �           u m     ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                   �#     ����x� H�]	    @�     J   J   ��     H�]	J                  2         �                 � � �           u m     ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                   �#     ����x� H�]	    @�     J   J   ��     H�]	J                  2         �                 � � �           u m     ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                   �#     ����x� H�]	    @�     J   J   ��     H�]	J                  2         �                 � � �           u m     ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                   �#     ����x� H�]	    @�     J   J   ��     H�]	J                  2         �                 � � �           u m     ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                   �#     ����x� H�]	    @�     J   J   ��     H�]	J                  2         �                 � � �           u m     ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                   �#     ����x� H�]	    @�     J   J   ��     H�]	J                  2         �                 � � �           u m     ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                   �#     ����x� H�]	    @�     J   J   ��     H�]	J                  2         �                 � � �           u m     ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                   �#     ����x� H�]	    @�     J   J   ��     H�]	J                  2         �                 � � �           u m     ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                   �#     ����x� H�]	    @�     J   J   ��     H�]	J                  2         �                 � � �           u m     ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                   �#     ����x� H�]	    @�     J   J   ��     H�]	J                  2         �                 � � �           u m     ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                   �#     ����x� H�]	    @�     J   J   ��     H�]	J                  2         �                 � � �           u m     ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                   �#     ����x� H�]	    @�     J   J   ��     H�]	J                  2         �                 � � �           u m     ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                               �� 	 CTitleBox        ��<    `�X                               �	                  �         �  @                  ���                                                  �  @  "�     <   �  <     ��                                                        "�     |   �  |     ��                                                       "�     �   �  �     ��    ���t                                                "�     �   �  �     ��                                                        8� h      t  4     ��                                                      h      t  4   h      t  4   [title]                                       8� �   H   �  x     ��                                                      �   H   �  x   �   H   �  x   [description]                                       8� P   �   X  �     ��                                                      P   �   X  �   P   �   X  �   [id]                                       8� �   �   �  �     ��                                                      �   �   �  �   �   �   �  �   
[designer]                                       8�      ]   1    ��        	                                                   ]   1       ]   1  Date :       ��  4  ��  �                  8� p     x  4   	 ��        
                                              p     x  4  p     x  4  [date]                                       8�       U   1    
 ��                                                            U   1         U   1   Title :       ��  4  ��  �                  8�    L   �   q     ��                                                         L   �   q      L   �   q   Description :       ��  �  ��  �                  8�    �   8   �     ��                                                         �   8   �      �   8   �   ID :       ��  �  8�  J                  8�    �   �   �     ��                                                         �   �   �      �   �   �   
Designer :       ��  t  p�  
                   LMNOPQRSTVWXYZ          U     	title box     Miscellaneous      �?    9 
 ��  CParamSubBehavior    
 ΁  ����        ��������΁  ����       ��������΁  ����       ��������΁  ����       ��������΁  ����       ��������΁  ����       ��������΁  ����       ��������΁  ����       ��������΁  ����       ��������΁  ����  	     ��������      
 9                      �               ������   CParamSubModelType�� ����  
   ��  	 CParmDefn            title                i�            description                i�            id                i�            designer                i�            Date :                i�            date                i�            Title :                i�            Description :                i�            ID :                i�            
Designer :                            ����             `         �?�� 	 CGraphDoc�  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                   H�����@{c�'�P�[����S@�W�UxO\����8S�
��o�             2         �                 � � �           ��    ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                         In1In2In3In4In5In6Out1Out2                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          1m  0                            100   100                                                           1m  0                            100   100                              1m  0                            100   100                              1m  0                            100   100                                                 
               1m  0                            100   100                            ��   CPartPackage     ��   CPackage�   DIP-14�14 pin dual in line package                                                                                                                                                                                                                               �     :;<=>?@ABCDEFGHI      ��   CMiniPartPin    ����ClrClr     INClr�  6@  z�   ����UpUp     INUp�  7@  z�   ����DownDown     INDown 	  8@  z�   ����LoadLoad     INLoad	  9@  z�   ����AA     INA	  :@  z�   ����BB     INB	  ;@  z�   ����CC     INC	  <@  z�   ����DD     IND	  =@  z�   ����COCO     OUTCO	  >@  z�	   ����BOBO     OUTBO	  ?@  z�
   ����QAQA     OUTQA	  @@  z�   ����QBQB     OUTQB		  A@  z�   ����QCQC     OUTQC
	  B@  z�   ����QDQD     OUTQD	  C@  74ALS192 (XSpice)74ALS192 (XSpice)��  CXSpiceBehavior       clrupdownloadabcdcoboqaqbqcqd ��   CBehPin 6@  clr����    �  clr����                         ���� 7@  up����   �  up����                         ���� 8@  down����   �  down����                         ���� 9@  load����   �  load����                         ���� :@  a����   �  a����                        ���� ;@  b����   �  b����                         ���� <@  c����   �  c����                         ���� =@  d����   �  d����                        ���� >@  co����   �  co����                        ���� ?@  bo����	   �  bo����                        ���� @@  qa����
   �  qa����                       ���� A@  qb����   �  qb����                        ���� B@  qc����   �  qc����                        ���� C@  qd����   �  qd����                       ��74192 ALS (XSpice)74192 ALS (XSpice)  8 X            ��������������Digital<   Generic                       * time value qaQAdownDownqbQBclrClrqcQCqdQDloadLoadupUpaAcoCObBboBOcCdD DdDowndownQAqaQBqbQCqcLoadloadQDqdClrclrUpupCOcoBOboAaBbCc                                                                                                                        z�    ����AA     INA  Q  InputInput                  z�    ����AA     INA  Q  InputInput                  z�    ����AA     INA  Q  InputInput                  z�    ����AA     INA  Q  InputInput                  z�    ����AA     INA  Q  InputInput                  z�    ����AA     INA  Q  InputInput               w z�    ����aA     IN1AA  �?  z�   ����bB     IN1BB  �?  z�   ����yY     OUT1Y@  �?     ��   CPackagePin 1 a   A1A�� 2 b   A1B�� 3 y   A1Y�� 4 a   B2A�� 5 b   B2B�� 6 y   B2Y�� 7  GND  COMGND�� 8 y   C3Y�� 9 a  	 C3A�� 10 b  
 C3B�� 11 y   D4Y�� 12 a   D4A�� 13 b   D4B�� 14  VCC  COMVCCXSpice 2input AND gateGatesGeneric=      7408 A74LS08NA1                        DIP1474LS08N74LS08N��       aby �� �?  a����    �  a����                        ���� �?  b����   �  b����                        ���� �?  y����   �  y����                        ��7408 LS 2-input And7408 LS 2-input And  8               ���Digital<   Generic                       * time value yYaAbB YyAaBb                                 Output_PortOutput_Port              z�    ����portport       ��������Output_PortOutput_Port                                                      l 