    � B2SPICE zzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzz      ��  CPart         @  `        @  `              74LS76N��  CIntPin    ��  CWire      �         �         @  `        @  `              74LS76N �   �    	 �   
   �
         @  `        @  `              74LS76N�          16 �   �    �        ��   TInPort       _   @         _   @                 Input ��  CExtPin    ��  CVertex   `   
   ��  CSegment?    �J      �
   �A   �K   �  �
   �@   �*   �  �   �   �   �  `   �    �U   �  `   �
   �   �  `   "     !                             �    �R      �   �J   �    �  �   &     %     $    
                                                @  �   A        `	          In3     ��   CPin                    ��                                                       �   @   A��  TEllipse �   8   �   H                  ����
[negative]               ���                    �   8   �   H   �   8   �   H   �� 
 TRectangle t       �   @                   ����A                                      t       �   @   ,� t   @   �   `                   ����A                                      t   @   �   `   ��  TLine �   @   �   @     ��                                                        ,�         �   `                   ����                                                 �   `   /� t       t   `     
 ��    ��W                                              ��  TPolygon                    ��                                                       ��  TPoint�   \    �  5��   P    @  5��   P    �  5��   D       5��   D        5��   P        5��   P    �}T    3�                    ��                                                       5��   $        5��   0    P��5��   0    �  5��   <    ��S5��   <    @  5��   0    �  5��   0    �|T    ��  
 TTextField �       �   8    	 ��        	                                               �       �   8   �       �   8   	[A.nbits]      <       ����            �      "Arial                �       �   8   E�    (      M     ��        
                                                 (      M      (      M   [value]       ,  �	  d  n
     (   l   P   E� ��������+   #     ��                                                       ��������+   #   ��������+   #   	[refname]         Q	  �  �	  ���������       ) 1   0   . =   G 4 F H -   + 2      input_general     Miscellaneous      �?      ��   TInPortModel       A ��  	 TModelPin Q  A����        A����                         ��             0��    ��������             0��    ��������             0��    ��������             0��    ��������             0��    ��������             0��    �������� d   :�0�yE>10e-9��    �������� d   :�0�yE>10e-9��    ��������                            ����  ����:�0�yE>10e-9��d         ����  ����:�0�yE>10e-9��d   �      J   �����         d   :�0�yE>10e-9��    �������� d   :�0�yE>10e-9��    ��������1 Bit Inport1 Bit Inport   �            L Digital<   Generic   In3In3           ����  ��    �������� ����  ��    �������� ����  ��    �������� ����  ��    �������� ����  ��    �������� ����  ��    �������� ����  ��    ��������          ����             In ��   CPartPin    ����AA      INAA�>      Digital Instruments Generic                         `   `              `   �  �              `   �   yE>       �  `   `          �      7 �        �         �  �        �  �              74LS04NO �   �
    �   R  
  10 Q  K� V  K����       K����                          ��      x��    ��������      x��    ��������      x��    ��������      x��    ��������      x��    ��������      x��    �������� d   :�0�yE>10e-9��    �������� d   :�0�yE>10e-9��    ��������                             ����  ����:�0�yE>10e-9��d         ����  ����:�0�yE>10e-9��d   �     R ��   TJKFFLS       SJClkKRQQ' K� S  S����        S����                          ��      x��    ��������      x��    ��������      x��    ��������      x��    ��������      x��    ��������      x��    �������� d   :�0�yE>10e-9��    �������� d   :�0�yE>10e-9��    ��������                            ����  ����:�0�yE>10e-9��d         ����  ����:�0�yE>10e-9��d   �      V   �����     ��   d   :�0�yE>10e-9��    �������� d   :�0�yE>10e-9��    ��������K� T  J����       J����                          ��      x��    ��������      x��    ��������      x��    ��������      x��    ��������      x��    ��������      x��    �������� d   :�0�yE>10e-9��    �������� d   :�0�yE>10e-9��    ��������                             ����  ����:�0�yE>10e-9��d         ����  ����:�0�yE>10e-9��d   �      V   �����     ��   d   :�0�yE>10e-9��    �������� d   :�0�yE>10e-9��    ��������K� U  Clk����       Clk����                          ��      x��    ��������      x��    ��������      x��    ��������      x��    ��������      x��    ��������      x��    �������� d   :�0�yE>10e-9��    �������� d   :�0�yE>10e-9��    ��������                           ����  ����:�0�yE>10e-9��d         ����  ����:�0�yE>10e-9��d   �     �    �   Z    11 �    Z    ��   TClock       �   �  �      �   �  �              Clock\ �    �9   �  @   �   �   `  @   a     `     �   ` �   �  @   �   d �%   �  �   �/   f �    �  �   g �   �#   �      �   j �Q          �I   �   �      m     l     k    
        i     h     �0   h �<    
  �   o �1   �:    
      q �-   r �)   �
      �C   �;   �      u     t     s                p     �   p �?   �  �   �4   �=   �      y �2   z �   @      �5   �I   �      }     |     {                x     w                         e         c                    �     A�                 U1     (�                   ��                                                       �   `   A,�     @   �   �                  ����                                             @   �   �   /� �   `   �   `     ��    �X                                                /� `   @   `   �     ��    8�W                                                /� p   h   x   h     ��    ��W                                                /� x   T   x   h     ��    X                                                /� x   T   �   T     ��    ��W                                                /� �   T   �   h     ��    �W                                                /� �   h   �   h     ��     X                                                /� �   P   �   p      ��    8�W	                                                E�    P   Z   u    
 ��        
                                                  P   Z   u      P   Z   u   [period]       P    0  �     P   P   t   E� �   `   �   �    	 ��                                                      �   `   �   �   �   `   �   �   ns          @  p  �  �   `   �   x   E�     �����        ��                                                           �����          �����      	[devname]        ����������������    �����      E�        *   @     ��                                                              *   @          *   @   	[refname]          h  �           �   <    �   �   �   �   � �   � � � �   �   �        �      Clock     Miscellaneous      �?      ��   TClockModel     ��  CValue �  I�����z>100n      ���������� �  I�����j>50n     �������� A K�     A����    ����A����                          ��      x��    ��������      x��    ��������      x��    ��������      x��    ��������      x��    ��������      x��    �������� d   :�0�yE>10e-9��    �������� d   :�0�yE>10e-9��    ��������                             ����  ����:�0�yE>10e-9��d         ����  ����:�0�yE>10e-9��d   �     Z �   �����         d   :�0�yE>10e-9��    �������� d   :�0�yE>10e-9��    ��������ClockClock              � Digital InstrumentsO   Generic   U1U1           ����  ��    �������� ����  ��    �������� ����  ��    �������� ����  ��    �������� ����  ��    �������� ����  ��    �������� ����  ��    ��������  al      ����Generic             U M�    ����AA      INAA�  ����Digital InstrumentsDigital Clock inputGeneric                                                                              �'                                   11 �   Z    11 �   Z    11  K� U  Clk����       Clk����                          ��      x��    ��������      x��    ��������      x��    ��������      x��    ��������      x��    ��������      x��    �������� d   :�0�yE>10e-9��    �������� d   :�0�yE>10e-9��    ��������                           ����  ����:�0�yE>10e-9��d         ����  ����:�0�yE>10e-9��d   �     Z U�       SJClkKRQQ' K� S  S����        S����                          ��      x��    ��������      x��    ��������      x��    ��������      x��    ��������      x��    ��������      x��    �������� d   :�0�yE>10e-9��    �������� d   :�0�yE>10e-9��    ��������                            ����  ����:�0�yE>10e-9��d         ����  ����:�0�yE>10e-9��d   �      �   �����     ��   d   :�0�yE>10e-9��    �������� d   :�0�yE>10e-9��    ��������K� T  J����       J����                          ��      x��    ��������      x��    ��������      x��    ��������      x��    ��������      x��    ��������      x��    �������� d   :�0�yE>10e-9��    �������� d   :�0�yE>10e-9��    ��������                             ����  ����:�0�yE>10e-9��d         ����  ����:�0�yE>10e-9��d   �     �    �   �    1 �   �    1 �    �    ��   TOutPort       _   @         _   @                 Output_Port� �    �   �   
   �'   �3   �   
   � �*   � �5   �  �   � �;   � �   �  �   � �8   �/   `  �   �     �                �3   � �$   @  �   �9   �N   �  �   �     �     �                        �     �(   � �4   �   
   �                        �   port     �  `	          Q1     (�                   ��                                                           @   port,�         �   `                   ����                                                 �   `   /�     @       @      ��                                                        *�    8       H                  ����
[negative]               ���                       8       H      8       H   E� (   ,   :   Q     ��                                                      (   ,   :   Q   (   ,   :   Q   [value]       X  �	  �  z
  (   ,   �   T   E�     $       <     ��                                                           $       <       $       <   [port.nbits]      <       ����            �      "Arial                    $       <   E�     ����M         ��                                                           ����M           ����M       	[refname]       @  H	  �  �	      �����       �   � � � � � �      Output_Port     Miscellaneous      �?      ��   TOutPortModel       port K� ����port����        port����                                         0��    ��������             0��    ��������             0��    ��������             0��    ��������             0��    ��������             0��    �������� d   :�0�yE>10e-9��    �������� d   :�0�yE>10e-9��    ��������                             ����  ����:�0�yE>10e-9��d         ����  ����:�0�yE>10e-9��d   �     � �   �����     ��   d   :�0�yE>10e-9��    �������� d   :�0�yE>10e-9��    ��������Output_PortOutput_Port   �            � Digital<   Generic   Q1Q1           ����  ��    �������� ����  ��    �������� ����  ��    �������� ����  ��    �������� ����  ��    �������� ����  ��    �������� ����  ��    ��������          ����       ����  Out M�    ����portport       A X]      Digital Instruments Generic                                                                                                             1  � � K� X  Q����       Q����                         �� �   :�0�yU>20ns��    ��������      x��    �������� �   ,i�)+P>15ns��    �������� �   :�0�yU>20ns��    ��������      x��    �������� �   ,i�)+P>15ns��    �������� d   :�0�yE>10e-9��    �������� d   :�0�yE>10e-9��    ��������                            ����  ����:�0�yE>10e-9��d         ����  ����:�0�yE>10e-9��d   �     � U�       SJClkKRQQ' K� S  S����        S����                          ��      x��    ��������      x��    ��������      x��    ��������      x��    ��������      x��    ��������      x��    �������� d   :�0�yE>10e-9��    �������� d   :�0�yE>10e-9��    ��������                            ����  ����:�0�yE>10e-9��d         ����  ����:�0�yE>10e-9��d   �      �   �����     ��   d   :�0�yE>10e-9��    �������� d   :�0�yE>10e-9��    ��������K� T  J����       J����                          ��      x��    ��������      x��    ��������      x��    ��������      x��    ��������      x��    ��������      x��    �������� d   :�0�yE>10e-9��    �������� d   :�0�yE>10e-9��    ��������                             ����  ����:�0�yE>10e-9��d         ����  ����:�0�yE>10e-9��d   �     
 �   �����     ��   d   :�0�yE>10e-9��    �������� d   :�0�yE>10e-9��    ��������K� U  Clk����       Clk����                          ��      x��    ��������      x��    ��������      x��    ��������      x��    ��������      x��    ��������      x��    �������� d   :�0�yE>10e-9��    �������� d   :�0�yE>10e-9��    ��������                           ����  ����:�0�yE>10e-9��d         ����  ����:�0�yE>10e-9��d   �     Z �   �����     ��   d   :�0�yE>10e-9��    �������� d   :�0�yE>10e-9��    ��������K� V  K����       K����                          ��      x��    ��������      x��    ��������      x��    ��������      x��    ��������      x��    ��������      x��    �������� d   :�0�yE>10e-9��    �������� d   :�0�yE>10e-9��    ��������                             ����  ����:�0�yE>10e-9��d         ����  ����:�0�yE>10e-9��d   �     �	    �   �  	  9 �   �  	  9  � K� Y  Q'����       Q'����                         �� �   :�0�yU>20ns��    ��������      x��    �������� �   ,i�)+P>15ns��    �������� �   :�0�yU>20ns��    ��������      x��    �������� �   ,i�)+P>15ns��    �������� d   :�0�yE>10e-9��    �������� d   :�0�yE>10e-9��    ��������                           ����  ����:�0�yE>10e-9��d         ����  ����:�0�yE>10e-9��d   �     � V   �����         d   :�0�yE>10e-9��    �������� d   :�0�yE>10e-9��    ��������	 9�   �����     ��   d   :�0�yE>10e-9��    �������� d   :�0�yE>10e-9��    ��������K� W  R����       R����                          ��      x��    ��������      x��    ��������      x��    ��������      x��    ��������      x��    ��������      x��    �������� d   :�0�yE>10e-9��    �������� d   :�0�yE>10e-9��    ��������                            ����  ����:�0�yE>10e-9��d         ����  ����:�0�yE>10e-9��d   �     �    �   �    12 �   �    12 �   �    12 �    �    �	       _   @         _   @                 Input� �    �   �
      �>   �G   `	      �     �     �=   � �B   @      �   �A   @  �   �   �"   @  �   � �F   � �O   @      � �6   �@   @  `   �     �        
            �     �     �     � �   � �H          �<   �C   �      �7   �D   �      � �)   � �   `      � �#   �E          �     �                    �     �     �     �   �!   �      �   � �0      `   �         �        �     �                    	        @  �   A   @  @          In1     (�                    ��                                                       �   @   A*� �   8   �   H                  ����
[negative]               ���                    �   8   �   H   �   8   �   H   ,� t       �   @                   ����A                                      t       �   @   ,� t   @   �   `                   ����A                                      t   @   �   `   /� �   @   �   @     ��                                                        ,�         �   `                   ����                                                 �   `   /� t       t   `     
 ��                                                      3�                    ��                                                       5��   \       5��   P       5��   P       5��   D       5��   D    `  5��   P       5��   P    `yW    3�                    ��                                                       5��   $       5��   0    `  5��   0        5��   <       5��   <    �  5��   0    �  5��   0    `xW    E� �       �   8    	 ��        	                                               �       �   8   �       �   8   	[A.nbits]      <       ����            �      "Arial                �       �   8   E�    (      M     ��        
                                                 (      M      (      M   [value]       L  �  �  N     (   l   P   E� ��������+   #     ��                                                       ��������+   #   ��������+   #   	[refname]       :  1  �  �  ���������       � �   �   � �    � � �   � �      input_general     Miscellaneous      �?      I�       A K�     A����    ����A����                         ��             0��    ��������             0��    ��������             0��    ��������             0��    ��������             0��    ��������             0��    �������� d   :�0�yE>10e-9��    �������� d   :�0�yE>10e-9��    ��������                            ����  ����:�0�yE>10e-9��d         ����  ����:�0�yE>10e-9��d   �     �   �����        d   :�0�yE>10e-9��    �������� d   :�0�yE>10e-9��    ��������1 Bit Inport1 Bit Inport   �t            Digital<   Generic   In1In1           ����  ��    �������� ����  ��    �������� ����  ��    �������� ����  ��    �������� ����  ��    �������� ����  ��    �������� ����  ��    ��������  Lo�    ����            In M�    ����AA      INAAQ  ����Digital Instruments Generic                         `   `              `   �  �              `   �             �  `   `          �      12  K� W  R����       R����                          ��      x��    ��������      x��    ��������      x��    ��������      x��    ��������      x��    ��������      x��    �������� d   :�0�yE>10e-9��    �������� d   :�0�yE>10e-9��    ��������                            ����  ����:�0�yE>10e-9��d         ����  ����:�0�yE>10e-9��d   �     � �   �����     ��   d   :�0�yE>10e-9��    �������� d   :�0�yE>10e-9��    ��������� K� W  R����       R����                          ��      x��    ��������      x��    ��������      x��    ��������      x��    ��������      x��    ��������      x��    �������� d   :�0�yE>10e-9��    �������� d   :�0�yE>10e-9��    ��������                            ����  ����:�0�yE>10e-9��d         ����  ����:�0�yE>10e-9��d   �     � V   �����     ��   d   :�0�yE>10e-9��    �������� d   :�0�yE>10e-9��    �������� 12�   �����     ��   d   :�0�yE>10e-9��    �������� d   :�0�yE>10e-9��    ��������� K� Y  Q'����       Q'����                         �� �   :�0�yU>20ns��    ��������      x��    �������� �   ,i�)+P>15ns��    �������� �   :�0�yU>20ns��    ��������      x��    �������� �   ,i�)+P>15ns��    �������� d   :�0�yE>10e-9��    �������� d   :�0�yE>10e-9��    ��������                           ����  ����:�0�yE>10e-9��d         ����  ����:�0�yE>10e-9��d   �     �    �      3 �      3  K� V  K����       K����                          ��      x��    ��������      x��    ��������      x��    ��������      x��    ��������      x��    ��������      x��    �������� d   :�0�yE>10e-9��    �������� d   :�0�yE>10e-9��    ��������                             ����  ����:�0�yE>10e-9��d         ����  ����:�0�yE>10e-9��d   �     �   �����     ��   d   :�0�yE>10e-9��    �������� d   :�0�yE>10e-9��    �������� 3�   �����         d   :�0�yE>10e-9��    �������� d   :�0�yE>10e-9��    ��������76/2 LS JK Neg Edge-Trig FF76/2 LS JK Neg Edge-Trig FF 0 [            � � � � � � Digital<   Analog Devices   A1A1           ���� x��    �������� ���� x��    �������� �'	 hUMu?60u��    �������� �r��b2U0*�C�-.6m��    �������� ���-C��6:�-.4m��    ��������  ������Mb�?8m��    ��������  Zb����Mbp?4m��    ��������          ����LS                 0��    �������� ����    8�|A30meg��    �������� �   vԷ1�X>23n��    �������� �   ����o�V>21n��    ��������  �����        d   :�0�yE>10e-9��    �������� d   :�0�yE>10e-9��    �������� 1�   �����     ��   d   :�0�yE>10e-9��    �������� d   :�0�yE>10e-9��    ��������� K� X  Q����       Q����                         �� �   :�0�yU>20ns��    ��������      x��    �������� �   ,i�)+P>15ns��    �������� �   :�0�yU>20ns��    ��������      x��    �������� �   ,i�)+P>15ns��    �������� d   :�0�yE>10e-9��    �������� d   :�0�yE>10e-9��    ��������                            ����  ����:�0�yE>10e-9��d         ����  ����:�0�yE>10e-9��d   �     �    �      5 �       ��       _   @         _   @                 Output_Port�    �   @   
   �%   �2   @  �	           �&   �   @  �   �$   �   �  �   �   �>   �  �                                             �   port     @  `	          Q0     (�                   ��                                                           @   port,�         �   `                   ����                                                 �   `   /�     @       @      ��                                                        *�    8       H                  ����
[negative]               ���                       8       H      8       H   E� (   ,   :   Q     ��                                                      (   ,   :   Q   (   ,   :   Q   [value]       �  �	  �  z
  (   ,   �   T   E�     $       <     ��                                                           $       <       $       <   [port.nbits]      <       ����            �      "Arial                    $       <   E�     ����M         ��                                                           ����M           ����M       	[refname]       �  H	  (  �	      �����          !     Output_Port     Miscellaneous      �?      ��       port K� ����port����        port����                                         0��    ��������             0��    ��������             0��    ��������             0��    ��������             0��    ��������             0��    �������� d   :�0�yE>10e-9��    �������� d   :�0�yE>10e-9��    ��������                             ����  ����:�0�yE>10e-9��d         ����  ����:�0�yE>10e-9��d   �     "  �����     ��   d   :�0�yE>10e-9��    �������� d   :�0�yE>10e-9��    ��������Output_PortOutput_Port   �            #Digital<   Generic   Q0Q0           ����  ��    �������� ����  ��    �������� ����  ��    �������� ����  ��    �������� ����  ��    �������� ����  ��    �������� ����  ��    ��������          ����       ����  Out M�    ����portport       A �>      Digital Instruments Generic                                                                                                             5  # 5�   �����        d   :�0�yE>10e-9��    �������� d   :�0�yE>10e-9��    ��������K� Y  Q'����       Q'����                         �� �   :�0�yU>20ns��    ��������      x��    �������� �   ,i�)+P>15ns��    �������� �   :�0�yU>20ns��    ��������      x��    �������� �   ,i�)+P>15ns��    �������� d   :�0�yE>10e-9��    �������� d   :�0�yE>10e-9��    ��������                           ����  ����:�0�yE>10e-9��d         ����  ����:�0�yE>10e-9��d   �     �    �   &   6  % 6�   �����         d   :�0�yE>10e-9��    �������� d   :�0�yE>10e-9��    ��������76/2 LS JK Neg Edge-Trig FF76/2 LS JK Neg Edge-Trig FF 0 [            � � � %Digital<   Analog Devices   A2A2           ���� x��    �������� ���� x��    �������� �'	 hUMu?60u��    �������� �r��b2U0*�C�-.6m��    �������� ���-C��6:�-.4m��    ��������  ������Mb�?8m��    ��������  Zb����Mbp?4m��    ��������          ����LS                 0��    �������� ����    8�|A30meg��    �������� �   vԷ1�X>23n��    �������� �   ����o�V>21n��    ��������  �����     ��   d   :�0�yE>10e-9��    �������� d   :�0�yE>10e-9��    ��������� � Y  11V   �����     ��   d   :�0�yE>10e-9��    �������� d   :�0�yE>10e-9��    ��������T K� X  Q����       Q����                         �� �   :�0�yU>20ns��    ��������      x��    �������� �   ,i�)+P>15ns��    �������� �   :�0�yU>20ns��    ��������      x��    �������� �   ,i�)+P>15ns��    �������� d   :�0�yE>10e-9��    �������� d   :�0�yE>10e-9��    ��������                            ����  ����:�0�yE>10e-9��d         ����  ����:�0�yE>10e-9��d   �     
 V   �����        d   :�0�yE>10e-9��    �������� d   :�0�yE>10e-9��    ��������� 76/2 LS JK Neg Edge-Trig FF76/2 LS JK Neg Edge-Trig FF 0 [            W X Y T (� Digital<   Analog Devices   A6A6           ���� x��    �������� ���� x��    �������� �'	 hUMu?60u��    �������� �r��b2U0*�C�-.6m��    �������� ���-C��6:�-.4m��    ��������  ������Mb�?8m��    ��������  Zb����Mbp?4m��    ��������          ����LS                 0��    �������� ����    8�|A30meg��    �������� �   vԷ1�X>23n��    �������� �   ����o�V>21n��    ��������  �����     ��   d   :�0�yE>10e-9��    �������� d   :�0�yE>10e-9��    ��������K� 8  Y����       Y����                         �� �   ,i�)+P>15ns��    ��������      x��    �������� d   :�0�yE>10ns��    �������� �   ,i�)+P>15ns��    ��������      x��    �������� Z   h�+e�SC>9ns��    �������� d   :�0�yE>10e-9��    �������� d   :�0�yE>10e-9��    ��������                           ����  ����:�0�yE>10e-9��d         ����  ����:�0�yE>10e-9��d   �     R ��   TAnd       InY K� 7  In����        In����                          ��      x��    ��������      x��    ��������      x��    ��������      x��    ��������      x��    ��������      x��    �������� d   :�0�yE>10e-9��    �������� d   :�0�yE>10e-9��    ��������                             ����  ����:�0�yE>10e-9��d         ����  ����:�0�yE>10e-9��d   �      +  �����     ��   d   :�0�yE>10e-9��    �������� d   :�0�yE>10e-9��    ��������)04/6 LS Inverter04/6 LS Inverter = �            ,)Digital<   Generic   A5A5           ���� x��    �������� ���� x��    �������� @ �h㈵��>20u��    �������� ���-C��6:�-.4m��    �������� ���-C��6:�-.4m��    ��������  ������Mb�?8m��    ��������  6nb2U0*�c?2.4m��    ��������          ����LS      �����        d   :�0�yE>10e-9��    �������� d   :�0�yE>10e-9��    ��������
 10 
 P 10 �    !        �  in    �   �X   `  `   �   �,      `   0 
   /    �   /�P      `   �G   �&   �  `   4 
   3    2 
  
         
        �  �  out    �  �
          A5     (�                   ��                                                           �   in(�                   ��                                                      �   �   out*� l   t   �   �                   ���                                          l   t   �   �   l   t   �   �   /� �   �   �   �     ��      �?                                                /�     �   ,   �     ��    �Cd                                                3� ����    ����      ��                                                         5�,   \    P��5�,   �        5�l   �        5�,   \    x�\    E� ����   �   0     ��                                                       ����   �   0   ����   �   0   	[devname]        ��������������������   �   0   E� ����0   >   X     ��                                                       ����0   >   X   ����0   >   X   	[refname]       t  p  <    ����0   �   T   	 8  6:7;@A9     Inverter    Inverter IEEEMiscellaneous      �?    =  +  A M�    ����inIn      INA1A�>      M�   ����outY      OUTA1Y�>     M�    ����inIn      INB1A�>      M�   ����outY      OUTB1Y�>     M�    ����inIn      INC1A�>      M�   ����outY      OUTC1Y�>     M�    ����inIn      IND1A����    M�   ����outY      OUTD1Y}	     M�    ����inIn      INE1A|	      M�   ����outY      OUTE1Y{	     M�    ����inIn      INF1Az	      M�   ����outY      OUTF1Y��W   Gatesdigital one-bit-wide inverterGenericDIP-14              7   L X , 7   7 � S �  � �    �T   @  �
   �   �
   @      �   �          �	   �W   �      �    U�   �  �
   V�   �'   `  �
   �   �      �
   Z     Y    X         W             T     S    �   S�      �
   �   �.   �  �
   ^         ]    \         R     Q    �"   �V          `         Q    P     O        
              S    �   %       �  J   �   l       @  Clk   �   3      �  K   �   �      `  R   �   �M   `	  �   �E   �8    
  �   �.   �6    
   
   �+   k�   �
   
   l�,   m�7   @   
   n                    j    i    �:   i�-   �
  �   �D   �F   @  �   r    q    p           h    g    �   �+   �  �   t    g       
      @  �  Q   �   �L   `	  `   �!   �    	  `   x 	   w    �   w�(   �
  `   �B   �1   @  `   | 	   {    z 	           	  
      @  �  Q'       �	          A6     (�                    ��                                                       `   `   S(�                   ��                                                          �   J(�                   ��                                                          �   Clk(�                   ��                                                          �   K(�                   ��                                                      `      R(�                   ��                                                      �   �   Q(�                   ��                                                      �   �   Q'/�     �   ,   �     ��    8�]                                                /� ,   �       �     ��    ����                                                ,�     �   �       	           	   ����                                             �   �      /�     �       �    
 ��    ����
                                                /�     �      �     ��    ����                                                /�     �       �     ��    ����                                                /� �   �   �   �     ��    `W�                                                /� �   �   �   �     ��                                                        *� X   p   h   �                  �                                           X   p   h   �   X   p   h   �   *� X      h                    �                                           X      h     X      h     /� `     `        ��    ����                                                *� �   �   �   �                  �                                           �   �   �   �   �   �   �   �   /� �   �   �   �     ��    �� �                                                *�    �       �                  �                                              �       �      �       �   /� `   `   `   p     ��    ����                                                E�    0   Z   X     ��                                                          0   Z   X      0   Z   X   	[refname]       h  P
  0  �
     0   �   T   E� (   �   0   �     ��                                                      (   �   0   �   (   �   0   �   j       �  p  �    (   �   p   �   E� 4   �   T   �     ��                                                      4   �   T   �   4   �   T   �   ck       �  �    f  4   �   |   �   E� (   �   8   �     ��                                                      (   �   8   �   (   �   8   �   k       �  0  �  �  (   �   p   �   E�       �   0     ��                                                             �   0         �   0   	[devname]        ����������������      �   0    ~���������������������      ����     7476 LS JK Neg Edge-Trig FF     7476 LS JK Neg Edge-Trig FF IEEEMiscellaneous      �?    0  V   A M�    ����SS      INAS�>      M�   ����JJ      INAJ�>     M�   ����ClkClk      INAClk�>     M�   ����KK      INAKh��   M�   ����RR      INAR�>     M�   ����QQ      OUTAQ�>     M�   ����Q'Q'      OUTAQ'�>     M�    ����SS      INBS�>      M�   ����JJ      INBJ�>     M�   ����ClkClk      INBClk�>     M�   ����KK      INBK����   M�   ����RR      INBR�>     M�   ����QQ      OUTBQ�>     M�   ����Q'Q'      OUTBQ'�>     
Flip Flops	flip flopGenericDIP-16              8 �    
    ��       _   @         _   @                 Output_Port��    m       �   port     �
  `	          Q2     (�                   ��                                                           @   port,�         �   `                   ����                                                 �   `   /�     @       @      ��                                                        *�    8       H                  ����
[negative]               ���                       8       H      8       H   E� (   ,   :   Q     ��                                                      (   ,   :   Q   (   ,   :   Q   [value]       �
  �	  0  z
  (   ,   �   T   E�     $       <     ��                                                           $       <       $       <   [port.nbits]      <       ����            �      "Arial                    $       <   E�     ����M         ��                                                           ����M           ����M       	[refname]       �
  H	  h  �	      �����       �  ������     Output_Port     Miscellaneous      �?      ��       port K� ����port����        port����                                         0��    ��������             0��    ��������             0��    ��������             0��    ��������             0��    ��������             0��    �������� d   :�0�yE>10e-9��    �������� d   :�0�yE>10e-9��    ��������                             ����  ����:�0�yE>10e-9��d         ����  ����:�0�yE>10e-9��d   �     
 �  �����     ��   d   :�0�yE>10e-9��    �������� d   :�0�yE>10e-9��    ��������Output_PortOutput_Port                 �Digital<   Generic   Q2Q2           ����  ��    �������� ����  ��    �������� ����  ��    �������� ����  ��    �������� ����  ��    �������� ����  ��    �������� ����  ��    ��������          ����       ����  Out M�    ����portport       A ����    Digital Instruments Generic                                                                                                             8  �� ( 8   8 � � � � 
�    _         S    �   q      �  J    �   t       @  Clk� l �   {      �  K��K�   �      `  R�����   �   @  �  Q 
  �   �   �  `   �   ��   @  `   �                    @  �  Q'�   �
  �	          A1     (�                    ��                                                       `   `   S(�                   ��                                                          �   J(�                   ��                                                          �   Clk(�                   ��                                                          �   K(�                   ��                                                      `      R(�                   ��                                                      �   �   Q(�                   ��                                                      �   �   Q'/�     �   ,   �     ��    ���                                                /� ,   �       �     ��    �K�                                                ,�     �   �       	           	   ����                                             �   �      /�     �       �    
 ��        
                                                /�     �      �     ��                                                        /�     �       �     ��    �dW                                                /� �   �   �   �     ��    JT                                                /� �   �   �   �     ��     �a                                                *� X   p   h   �                  �                                           X   p   h   �   X   p   h   �   *� X      h                    �                                           X      h     X      h     /� `     `        ��    8�\                                                *� �   �   �   �                  �                                           �   �   �   �   �   �   �   �   /� �   �   �   �     ��    (��                                                *�    �       �                  �                                              �       �      �       �   /� `   `   `   p     ��    �U                                                E�    0   Z   X     ��                                                          0   Z   X      0   Z   X   	[refname]       �
  P
  �  �
     0   �   T   E� (   �   0   �     ��                                                      (   �   0   �   (   �   0   �   j       �
  p      (   �   p   �   E� 4   �   T   �     ��                                                      4   �   T   �   4   �   T   �   ck         �  |  f  4   �   |   �   E� (   �   8   �     ��                                                      (   �   8   �   (   �   8   �   k       �
  0  (  �  (   �   p   �   E�       �   0     ��                                                             �   0         �   0   	[devname]        ����������������      �   0    �����������������������      ����     7476 LS JK Neg Edge-Trig FF     7476 LS JK Neg Edge-Trig FF IEEEMiscellaneous      �?    0  �   A M�    ����SS      INAS�>      M�   ����JJ      INAJ�>     M�   ����ClkClk      INAClkx��   M�   ����KK      INAKyE>   M�   ����RR      INAR ���   M�   ����QQ      OUTAQ d    M�   ����Q'Q'      OUTAQ'      M�    ����SS      INBS J�    M�   ����JJ      INBJ10e-   M�   ����ClkClk      INBClk0e-9   M�   ����KK      INBK  x   M�   ����RR      INBR      M�   ����QQ      OUTBQ 5   M�   ����Q'Q'      OUTBQ'      
Flip Flops	flip flopGenericDIP-16             16 �         �       _   @         _   @                 Input��    a   @  �   A (A �  `          In4     (�                    ��                                                       �   @   A*� �   8   �   H                  ����
[negative]               ���                    �   8   �   H   �   8   �   H   ,� t       �   @                   ����A                                      t       �   @   ,� t   @   �   `                   ����A                                      t   @   �   `   /� �   @   �   @     ��                                                        ,�         �   `                   ����                                                 �   `   /� t       t   `     
 ��                                                      3�                    ��                                                       5��   \    �  5��   P    @  5��   P    �  5��   D       5��   D        5��   P        5��   P    �}T    3�                    ��                                                       5��   $        5��   0    P��5��   0    �  5��   <    ��S5��   <    @  5��   0    �  5��   0    �|T    E� �       �   8    	 ��        	                                               �       �   8   �       �   8   	[A.nbits]      <       ����            �      "Arial                �       �   8   E�    (      M     ��        
                                                 (      M      (      M   [value]       �  �    n     (   l   P   E� ��������+   #     ��                                                       ��������+   #   ��������+   #   	[refname]       �  Q  B  �  ���������       ��  �  ��  ��  ��     input_general     Miscellaneous      �?      I�       A K� Q  A����        A����                         ��             0��    ��������             0��    ��������             0��    ��������             0��    ��������             0��    ��������             0��    �������� d   :�0�yE>10e-9��    �������� d   :�0�yE>10e-9��    ��������                            ����  ����:�0�yE>10e-9��d         ����  ����:�0�yE>10e-9��d   �        �����         d   :�0�yE>10e-9��    �������� d   :�0�yE>10e-9��    ��������1 Bit Inport1 Bit Inport   �            Digital<   Generic   In4In4           ����  ��    �������� ����  ��    �������� ����  ��    �������� ����  ��    �������� ����  ��    �������� ����  ��    �������� ����  ��    ��������  al      ����             In M�    ����AA      INAA����    Digital Instruments Generic                         `   `              `   �  �              `   �   yE>       �  `   `          �      16   � � W   16  �� 16 � [ 	� '�    Y         S> l �   �       �  J   �   |       @  Clk_�K�   �      �  K�����   �      `  R~R�K�     @  �  Q�����   �	   �  `   �H   �S   �  `                    @  �  Q'     @  �	          A2     (�                    ��                                                       `   `   S(�                   ��                                                          �   J(�                   ��                                                          �   Clk(�                   ��                                                          �   K(�                   ��                                                      `      R(�                   ��                                                      �   �   Q(�                   ��                                                      �   �   Q'/�     �   ,   �     ��                                                        /� ,   �       �     ��                                                        ,�     �   �       	           	   ����                                             �   �      /�     �       �    
 ��    ���t
                                                /�     �      �     ��    
                                                  /�     �       �     ��                                                        /� �   �   �   �     ��    �                                                  /� �   �   �   �     ��                                                        *� X   p   h   �                  �                                           X   p   h   �   X   p   h   �   *� X      h                    �                                           X      h     X      h     /� `     `        ��                                                        *� �   �   �   �                  �                                           �   �   �   �   �   �   �   �   /� �   �   �   �     ��                                                       *�    �       �                  �                                              �       �      �       �   /� `   `   `   p     ��                                                        E�    0   Z   X     ��                                                          0   Z   X      0   Z   X   	[refname]       �  P
  P  �
     0   �   T   E� (   �   0   �     ��                                                      (   �   0   �   (   �   0   �   j       �  p  �    (   �   p   �   E� 4   �   T   �     ��                                                      4   �   T   �   4   �   T   �   ck       �  �  <  f  4   �   |   �   E� (   �   8   �     ��                                                      (   �   8   �   (   �   8   �   k       �  0  �  �  (   �   p   �   E�       �   0     ��                                                             �   0         �   0   	[devname]        ����������������      �   0     !"#$()*      +%&'     7476 LS JK Neg Edge-Trig FF     7476 LS JK Neg Edge-Trig FF IEEEMiscellaneous      �?    0  �   A M�    ����SS      INAS�>      M�   ����JJ      INAJ�>     M�   ����ClkClk      INAClk��   M�   ����KK      INAK~A     M�   ����RR      INAR�>     M�   ����QQ      OUTAQ       M�   ����Q'Q'      OUTAQ'�>     M�    ����SS      INBS�>      M�   ����JJ      INBJ�>     M�   ����ClkClk      INBClk����   M�   ����KK      INBK�>     M�   ����RR      INBR   �   M�   ����QQ      OUTBQ�<�   M�   ����Q'Q'      OUTBQ'       
Flip Flops	flip flopGenericDIP-16                 ^ ��  �    �P     � Z � & 
 � R K H K       P$ ��   �            :    �   �       :        R\T"   �  � � i w ^k c 2a � XZe 0� tzVx`� � � � � lns jg o q { � y } � � � � p� � � �    |u rh� 4m & Y T Y h n   ;<        QSb � �y][� | �# � m� W d  ' � � j � f 5Y{t  u1q_� � }� � � koi` r v p z x � � � � � � s� � ~   wg� � 3l % O! aU/             
 ��@ ����        ����������             0     ���������� ����      @5     ����������  ʚ;�������?.1     ����������@ ����       ���������� ����       ���������� ����       ���������� ����       ���������� ���� true
     ���������� ����  false     ��������               
                  �� ����        ���������� ����       ����������  ����       ����������@ ����       ����������@ ����       ��������               
                  �� ����        ���������� ����       ����������@ ����       ����������  ����       ���������� ����       ���������� ����       ���������� ����       ���������� ����       ���������� ����       ���������� ����       ���������� ����       ��������               
                 �� ����dec     ���������� ����     @�@1k     ���������� ����    ��.A1meg     ���������� ����       20     ���������� ���� true     ���������� ���� true     ���������� ���� true	     ���������� ����  false
     ��������               
                 ��  ����        ����������  ����       ����������  ����       ���������� ����dec     ���������� ����       ���������� ����       ���������� ����  	     ���������� ����  
     ��������               
                  	 �� ����        ���������� ����       ���������� ����       ���������� ����       ���������� ����       ���������� ����       ���������� ����       ���������� ����       ���������� ����       ��������               
                 �� ����        ���������� ����       ���������� ����       ���������� ����dec     ���������� ����       ��������               
                     ��             0      ���������� ��� ����MbP?1m     ���������� �� �h㈵��>10u     ���������� '  ���ư>1u     ���������� ���� true     ���������� ����  false     ���������� ���� true     ���������� ����  false     ��������               
                 �� ����     @�@1K      ����������  ����       ����������  ����       ����������  ����       ��������               
         ��              ��  ����        ��������              
                  ��  ����        ��������              
                                  
                 ��@ ����        ����������@ ����       ���������� ����       ���������� ����       ���������� ����       ���������� ����       ���������� ����       ���������� ����       ���������� ����       ���������� ���� true	     ���������� ����  false
     ���������� ���� true     ���������� ����  false     ��������               
                 �� ����       5      ���������� ����       5     ���������� ����       5     ���������� ����       5     ���������� ����       ���������� ����  	     ���������� ����  
     ���������� ����       ���������� ����       ���������� ����       ���������� ���� true     ����������@ ����       ����������@ ����       ���������� ����       ���������� ����       ���������� ����       ���������� ����dec     ���������� ����       ���������� ����       ���������� ����       ���������� ���� true     ���������� ���� true     ���������� ���� true     ���������� ����  false     ���������� ���� true     ���������� ����  false      ���������� ���� true!     ���������� ����  false"     ��������               
                        �� ����       5      ���������� ����       5     ���������� ����       5     ���������� ����       5     ���������� ����       ���������� ����  	     ���������� ����  
     ���������� ����       ���������� ����       ���������� ����       ���������� ���� true     ����������@ ����       ����������@ ����       ���������� ����       ���������� ����       ���������� ����       ���������� ����dec     ���������� ����       ���������� ����       ���������� ����       ���������� ���� true     ���������� ���� true     ���������� ���� true     ���������� ����  false     ���������� ���� true     ���������� ����  false      ���������� ���� true!     ���������� ����  false"     ��������               
                 �� ����       5      ���������� ����       5     ���������� ����       5     ���������� ����       5     ���������� ����       ���������� ����  	     ���������� ����  
     ���������� ����       ���������� ����       ���������� ����       ���������� ���� true     ����������@ ����       ����������@ ����       ���������� ����       ���������� ����       ���������� ����       ���������� ����dec     ���������� ����       ���������� ����       ���������� ����       ���������� ���� true     ���������� ���� true     ���������� ���� true     ���������� ����  false     ���������� ���� true     ���������� ����  false      ���������� ���� true!     ���������� ����  false"     ��������               
                 �� ����       5      ���������� ����       5     ���������� ����       5     ���������� ����       5     ���������� ����       ���������� ����  	     ���������� ����  
     ���������� ����       ���������� ����       ���������� ����       ���������� ���� true     ����������@ ����       ����������@ ����       ���������� ����       ���������� ����       ���������� ����       ���������� ����dec     ���������� ����       ���������� ����       ���������� ����       ���������� ���� true     ���������� ���� true     ���������� ���� true     ���������� ����  false     ���������� ���� true     ���������� ����  false      ���������� ���� true!     ���������� ����  false"     ��������               
                 ��@ ����        ����������@ ����       ���������� ����       ���������� ����       ���������� ����       ���������� ����       ���������� ����       ���������� ����       ���������� ����decade     ���������� ���� true     ���������� ���� true     ���������� ���� true     ���������� ����  false     ��������               
                 �� ����        ���������� ����       ����������@ ����       ����������  ����       ���������� ����       ���������� ����       ���������� ����       ���������� ����       ���������� ����       ���������� ����       ���������� ����       ��������               
                        �� ����dec     ���������� ����     @�@1k     ���������� ����    ��.A1meg     ���������� ����       20     ���������� ����        0     ���������� ����        0     ���������� ���� true	     ���������� ���� true
     ���������� ����      I@50     ���������� ���� true     ���������� ����  false     ��������               
                          / �� ���� x'     ����������     �-���q=1E-12     ���������� @B -C��6?1E-4     ���������� ���� x     ���������� ���� x     ���������� ���� x     ���������� ���� x     ���������� ���� x     ���������� ���� x     ���������� ���� x	     ���������� ���� x!     ���������� ����    �  500
     ���������� ���� x     ���������� ����    �  500     ���������� ���� x$     ���������� ���� x$     ���������� ���� x%     ���������� ���� x"     ����������  ���� x*     ���������� ���� x     ���������� ���� x     ���������� ���� x     ���������� ���� x&     ���������� ���� x     ���������� ���� x     ���������� ���� x     ���������� ���� x+     ���������� ���� x,     ���������� ���� x-     ���������� ���� xg     ���������� ���� xf     ���������� ���� xd     ���������� ���� xe     ���������� ���� xh     ���������� ���� xj     ���������� ���� xi     ���������� ���� xk     ���������� ����    e��A1Gl     ����������             0�     ���������� ����      @5�     ���������� ����      @2.5�     ���������� ����      �?.5�     ���������� ����      @4.5�     ���������� 
   ��&�.>1n�     ���������� 
   ��&�.>1n�     ���������� 
   ��&�.>1n�     ���������� 
   ��&�.>1n�     ��������                                  Ariald        �ڬtĢ�h�  ۬t� ���t    �ڬtĢ�h�  ۬t� ���t ��  COpAnal                         
                        ����                                   �ڬtĢ�h�  ۬t� ���t    �ڬtĢ�h�  ۬t� ���t ��  CDCsweep       
 =>?@ABCDEF               
                      ����                                   �ڬtĢ�h�  ۬t� ���t    �ڬtĢ�h�  ۬t� ���t ��  CACsweep        WXYZ[\]^               
                      ����                                  �ڬtĢ�h�  ۬t� ���t    �ڬtĢ�h�  ۬t� ���t �� 
 CTranSweep        uvwxyz{|               
                      ����                                   �ڬtĢ�h�  ۬t� ���t    �ڬtĢ�h�  ۬t� ���t ��  CACdisto        pqrst               
                          ����                                  �ڬtĢ�h�  ۬t� ���t    �ڬtĢ�h�  ۬t� ���t Z�        �� ����        ���������� ����       ���������� ����       ���������� ����dec     ���������� ����       ��������               
         �                ����                                  �ڬtĢ�h�  ۬t� ���t    �ڬtĢ�h�  ۬t� ���t Z�        �� ����        ���������� ����       ���������� ����       ���������� ����dec     ���������� ����       ��������               
                         ����                                  �ڬtĢ�h�  ۬t� ���t    �ڬtĢ�h�  ۬t� ���t Z�        �� ����        ���������� ����       ���������� ����       ���������� ����dec     ���������� ����       ��������               
                          ����                                  �ڬtĢ�h�  ۬t� ���t    �ڬtĢ�h�  ۬t� ���t Z�        �� ����        ���������� ����       ���������� ����       ���������� ����dec     ���������� ����       ��������               
         �                ����                                  �ڬtĢ�h�  ۬t� ���t    �ڬtĢ�h�  ۬t� ���t Z�        �� ����        ���������� ����       ���������� ����       ���������� ����dec     ���������� ����       ��������               
                     	    ����                                  �ڬtĢ�h�  ۬t� ���t    �ڬtĢ�h�  ۬t� ���t ��  CACnoise        _`abcdef               
                   
    ����                                  �ڬtĢ�h�  ۬t� ���t    �ڬtĢ�h�  ۬t� ���t z�         ��  ����        ����������  ����       ����������  ����       ���������� ����dec     ���������� ����       ���������� ����       ���������� ����  	     ���������� ����  
     ��������              
                        ����                                  �ڬtĢ�h�  ۬t� ���t    �ڬtĢ�h�  ۬t� ���t ��  CFourier        }~�               
         ��                  ����                                   �ڬtĢ�h�  ۬t� ���t    �ڬtĢ�h�  ۬t� ���t ��  CACpz        	 ghijklmno               
                       ����                                   �ڬtĢ�h�  ۬t� ���t    �ڬtĢ�h�  ۬t� ���t ��  CDCtf         GHIJK               
                       ����                                   �ڬtĢ�h�  ۬t� ���t    �ڬtĢ�h�  ۬t� ���t ��  CDCsens         LMNOPQRSTUV               
                       ����                                   �ڬtĢ�h�  ۬t� ���t    �ڬtĢ�h�  ۬t� ���t                 ����                                   �ڬtĢ�h�  ۬t� ���t    �ڬtĢ�h�  ۬t� ���t ��  CShow         �              
                       ����                                   �ڬtĢ�h�  ۬t� ���t    �ڬtĢ�h�  ۬t� ���t ��  CShowmod         �              
                       ����                                   �ڬtĢ�h�  ۬t� ���t    �ڬtĢ�h�  ۬t� ���t �� 
 CLinearize        ��  ����        ��������               
                      ����                                   �ڬtĢ�h�  ۬t� ���t    �ڬtĢ�h�  ۬t� ���t ��  CParamTranSweep        �������������               
                      ����                                   �ڬtĢ�h�  ۬t� ���t    �ڬtĢ�h�  ۬t� ���t U             ����                                   �ڬtĢ�h�  ۬t� ���t    �ڬtĢ�h�  ۬t� ���t ��  CParamACSweep         	
               
                      ����                                  �ڬtĢ�h�  ۬t� ���t    �ڬtĢ�h�  ۬t� ���t ��  CMonteCarlo_op        ����������������������������               
                             ����                                   �ڬtĢ�h�  ۬t� ���t    �ڬtĢ�h�  ۬t� ���t ��  CMonteCarlo_dc        ����������������������������               
                      ����                                   �ڬtĢ�h�  ۬t� ���t    �ڬtĢ�h�  ۬t� ���t ��  CMonteCarlo_ac        ����������������������������               
                      ����                                  �ڬtĢ�h�  ۬t� ���t    �ڬtĢ�h�  ۬t� ���t ��  CMonteCarlo_tran        ����������������������������               
                      ����                                   �ڬtĢ�h�  ۬t� ���t    �ڬtĢ�h�  ۬t� ���t ��  CACsens                       
                             ����                                  �ڬtĢ�h�  ۬t� ���t    �ڬtĢ�h�  ۬t� ���t ��  CNetworkAnalysis         !"               
                      ����                                  �ڬtĢ�h�  ۬t� ���t    �ڬtĢ�h�  ۬t� ���t                 ����                                 >           ��   CDigSimResTemplate                     ��   TDigitalSignal            U1    ���� ����                        ��            Q2    ���� ����                        ��            Q1    ���� ����                        ��            Q0    ���� ����                        ��            In1    ���� ����                        ��            In3    ���� ����                        ��            In4    ���� ����                                  ���       ����  ����:�0�yU>+20.00n���   ����                       Arial����                       Arial����                       Arial                                          ����  ����        0��          ����  ����        0��                     �               ����  �����      1000������          0.000000e+000��    ��������      0.000000e+000��    ��������      0.000000e+000��    ��������   ����                       Arial����                       Arial����                       Arial����                       Arial                        �     �   �  �                     ����  ��    ��������   �   DIP-16�16 pin DIP                                                                                                                                                                                                                                                �     ��   CPackageAliasSuperPCBStandardDIP16      ��EagleBURR.LBRDIP-16      ��Orcad DIP.100/16/W.300/L.800      ��Pads DIP16      ��	UltiboardUltilib.l55DIP16      ��Eagleburr-brown.lbrDIL16      ��Eagledil.lbrDIL16     ��Eagle74xx-usDIL16      ��Eagle	74ttl-dinDIL16      ��EaglemaximDIL16      ��EagleeclDIL16      ��EagleexarDIL16      ��EaglefifoDIL16      ��Eagle
ic-packageDIL16      ��EaglelinearDIL16      ��EaglememoryDIL16      ��Eaglememory-hitachiDIL16      ��Eagle
memory-idtDIL16      ��Eagle
memory-necDIL16      ��Eaglemicro-harrisDIL16      ��Eaglemicro-intelDIL16      ��Eaglemicro-motorolaDIL16      ��Eaglemicro-philipsDIL16      ��EagleoptocouplerDIL16      ��Eagleopto-micro-linearDIL16      ��EagletexasDIL16      ��Eagleresistor-dilDIL16      ��Eaglest-microelectronicsDIL16      ��Eagletransistor-npnDIL16      ��Eagleuln-udnDIL16      ��Eagle
74ac-logicDIL16              A                                                                            �   DIP-16�16 pin DIP                                                                                                                                                                                                                                                �     �������������������������������        B                            �   DIP-16�16 pin DIP                                                                                                                                                                                                                                                �     �������������������������������        A                            �   DIP-14�14 pin dual in line package                                                                                                                                                                                                                               �     ��SuperPCBStandardDIP14      ��EagleBURR.LBRDIP-14      ��Orcad DIP.100/14/W.300/L.700      ��Pads DIP14      ��	UltiboardUltilib.l55DIP14      ��Eagleburr-brown.lbrDIL14      ��Eagledil.lbrDIL14     ��Eagleanalog-devicesDIL14      ��Eagle74xx-usDIL14      ��Eagle	74ttl-dinDIL14      ��EaglemaximDIL14      ��EagleexarDIL14      ��Eagle
ic-packageDIL14      ��Eagleresistor-dilDIL14      ��EagletexasDIL14      ��Eagle
74ac-logicDIL14              A    �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                   �#     ����d� ��_	    ,�     N   N   z�     ��_	N                  2         �                 � � �           u m     ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                   �#     ����d� ��_	    ,�     N   N   z�     ��_	N                  2         �                 � � �           u m     ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                   �#     ����d� ��_	    ,�     N   N   z�     ��_	N                  2         �                 � � �           u m     ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                   �#     ����d� ��_	    ,�     N   N   z�     ��_	N                  2         �                 � � �           u m     ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                   �#     ����d� ��_	    ,�     N   N   z�     ��_	N                  2         �                 � � �           u m     ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                   �#     ����d� ��_	    ,�     N   N   z�     ��_	N                  2         �                 � � �           u m     ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                   �#     ����d� ��_	    ,�     N   N   z�     ��_	N                  2         �                 � � �           u m     ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                   �#     ����d� ��_	    ,�     N   N   z�     ��_	N                  2         �                 � � �           u m     ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                   �#     ����d� ��_	    ,�     N   N   z�     ��_	N                  2         �                 � � �           u m     ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                   �#     ����d� ��_	    ,�     N   N   z�     ��_	N                  2         �                 � � �           u m     ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                   �#     ����d� ��_	    ,�     N   N   z�     ��_	N                  2         �                 � � �           u m     ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                   �#     ����d� ��_	    ,�     N   N   z�     ��_	N                  2         �                 � � �           u m     ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                   �#     ����d� ��_	    ,�     N   N   z�     ��_	N                  2         �                 � � �           u m     ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                   �#     ����d� ��_	    ,�     N   N   z�     ��_	N                  2         �                 � � �           u m     ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                   �#     ����d� ��_	    ,�     N   N   z�     ��_	N                  2         �                 � � �           u m     ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                   �#     ����d� ��_	    ,�     N   N   z�     ��_	N                  2         �                 � � �           u m     ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                   �#     ����d� ��_	    ,�     N   N   z�     ��_	N                  2         �                 � � �           u m     ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                   �#     ����d� ��_	    ,�     N   N   z�     ��_	N                  2         �                 � � �           u m     ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                   �#     ����d� ��_	    ,�     N   N   z�     ��_	N                  2         �                 � � �           u m     ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                   �#     ����d� ��_	    ,�     N   N   z�     ��_	N                  2         �                 � � �           u m     ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                   �#     ����d� ��_	    ,�     N   N   z�     ��_	N                  2         �                 � � �           u m     ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                   �#     ����d� ��_	    ,�     N   N   z�     ��_	N                  2         �                 � � �           u m     ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                   �#     ����d� ��_	    ,�     N   N   z�     ��_	N                  2         �                 � � �           u m     ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                   �#     ����d� ��_	    ,�     N   N   z�     ��_	N                  2         �                 � � �           u m     ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                   �#     ����d� ��_	    ,�     N   N   z�     ��_	N                  2         �                 � � �           u m     ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                   �#     ����d� ��_	    ,�     N   N   z�     ��_	N                  2         �                 � � �           u m     ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                   �#     ����d� ��_	    ,�     N   N   z�     ��_	N                  2         �                 � � �           u m     ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                   �#     ����d� ��_	    ,�     N   N   z�     ��_	N                  2         �                 � � �           u m     ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                   �#     ����d� ��_	    ,�     N   N   z�     ��_	N                  2         �                 � � �           u m     ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                   �#     ����d� ��_	    ,�     N   N   z�     ��_	N                  2         �                 � � �           u m     ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                               �� 	 CTitleBox                                                      �	                  ,�         �  @                  ���                                                  �  @  /�     <   �  <     ��                                                        /�     |   �  |     ��                                                        /�     �   �  �     ��    � <                                                 /�     �   �  �     ��                                                        E� h      t  4     ��                                                      h      t  4   h      t  4   [title]                                       E� �   H   �  x     ��                                                      �   H   �  x   �   H   �  x   [description]                                       E� P   �   X  �     ��                                                      P   �   X  �   P   �   X  �   [id]                                       E� �   �   �  �     ��                                                      �   �   �  �   �   �   �  �   
[designer]                                       E�      ]   1    ��        	                                                   ]   1       ]   1  Date :       �	  4  �
  �                  E� p     x  4   	 ��        
                                              p     x  4  p     x  4  [date]                                       E�       U   1    
 ��                                                            U   1         U   1   Title :       �	  4  �
  �                  E�    L   �   q     ��                                                         L   �   q      L   �   q   Description :       �	  �  �  �                  E�    �   8   �     ��                                                         �   8   �      �   8   �   ID :       �	  �  8
  J                  E�    �   �   �     ��                                                         �   �   �      �   �   �   
Designer :       �	  t  p  
                   ��������������          �     	title box     Miscellaneous      �?    9 
 ��  CParamSubBehavior    
 ��  ����        ����������  ����       ����������  ����       ����������  ����       ����������  ����       ����������  ����       ����������  ����       ����������  ����       ����������  ����       ����������  ����  	     ��������        9                                      ������   CParamSubModelType�� ����  
   ��  	 CParmDefn            title                ��            description                ��            id                ��            designer                ��            Date :                ��            date                ��            Title :                ��            Description :                ��            ID :                ��            
Designer :                            ����             `         �?�� 	 CGraphDoc�  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                                                                                            2         �                 � � �                   ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                         U1Q2Q1Q0In1In3In4                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              1m  0                            100   100                                                           1m  0                            100   100                              1m  0                            100   100                              1m  0                            100   100                                                 
               1m  0                            100   100                            ��   CPartPackage   ��   CPackage�   DIP-14�14 pin dual in line package                                                                                                                                                                                                                               �     ����������������   
��    ��   DIP-16�16 pin DIP                                                                                                                                                                                                                                                �     �������������������������������   
��        ��   CMiniPartPin    ����SS     INS�      �   ����JJ     INJ�     �   ����ClkClk     INClk�     �   ����KK     INK�     �   ����RR     INR�     �   ����QQ     OUTQ�     �   ����Q'Q'     OUTQ'�         ��   CPackagePin 4 J   A1J� 12 K   B2K� 1 Clk   A1CLK� 2 S   A~1PR� 3 R   A~1CLR� 11 Q   B2Q� 10 Q'  
 B~2Q� 5  VCC  COMVCC� 6 Clk   B2CLK� 7 S   B~2PR� 8 R   B~2CLR� 9 J  	 B2J� 13  GND  COMGND� 14 Q'   A~1Q� 15 Q   A1Q� 16 K   A1K	flip flop
Flip FlopsGenericC      7476 A74LS76NA1                DIP1674LS76N74LS76N                                                                  �    ����AA     INA  Q  InputInput                  �    ����AA     INA�      ClockClock                  �    ����portport       ��������Output_PortOutput_Port                  �    ����portport       ��������Output_PortOutput_Port                  �    ����portport       ��������Output_PortOutput_Port                �    ����SS     INS�      �   ����JJ     INJ�     �   ����ClkClk     INClk�     �   ����KK     INK�     �   ����RR     INR�     �   ����QQ     OUTQ�     �   ����Q'Q'     OUTQ'�          � 4 J   A1J� 12 K   B2K� 1 Clk   A1CLK� 2 S   A~1PR� 3 R   A~1CLR� 11 Q   B2Q� 10 Q'  
 B~2Q� 5  VCC  COMVCC� 6 Clk   B2CLK� 7 S   B~2PR� 8 R   B~2CLR� 9 J  	 B2J� 13  GND  COMGND� 14 Q'   A~1Q� 15 Q   A1Q� 16 K   A1K	flip flop
Flip FlopsGenericC      7476 A74LS76NA5               DIP1674LS76N74LS76N                                                                  �    ����AA     INA      InputInput                �    ����SS     INS�      �   ����JJ     INJ�     �   ����ClkClk     INClk�     �   ����KK     INK�     �   ����RR     INR�     �   ����QQ     OUTQ�     �   ����Q'Q'     OUTQ'�          6789:;<=>?@ABCDE	flip flop
Flip FlopsGenericC      7476 A74LS76NA5               DIP1674LS76N74LS76N��  CXSpiceBehavior       jkclksetresetoutNout ��   CBehPin }A  j����    �  j����                         ��P� ~A  k����   �  k����                         ��P� A  clk����   �  clk����                         ��P� "E  set����   �  set����                         ��P� �A  reset����   �  reset����                         ��P� �A  out����   �  out����                        ��P� �A  Nout����   �  Nout����                        ��7476 LS (Xspice)7476 LS (Xspice)  8 �t            QRSTUVWDigital<   Generic                       * time value jJkKresetRoutQsetSclkClkNoutQ' JjKkQ'NoutQoutRresetClkclkSset                                                                �    ����AA     INA  Q  InputInput                �    ����inIn     IN1A�  �>  �   ����outY     OUT1Y�  �>   P   � 1 in   A1A� 2 out   A1Y� 3 in   B2A� 4 out   B2Y� 5 in   C3A� 6 out   C3Y� 7  GND  COMGND� 8 out   D4Y� 9 in  	 D4A� 10 out  
 E5Y� 11 in   E5A� 12 out   F6Y� 13 in   F6A� 14  VCC  COMVCCdigital one-bit-wide inverterGatesGeneric=      7404 A74LS04NA4                                DIP1474LS04N74LS04NN�       inout P� �>  in����    �  in����                         ��P� �>  out����   �  out����                        ��7404 LS Inverter7404 LS Inverter  8               jkDigital<   Generic                       * time value inInoutY IninYout                                                               